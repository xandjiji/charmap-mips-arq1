module font_ROM(
    input wire dclk,                // clock (nao tenho certeza se eh esse que devo usar)
    input wire [10:0] char_select,  // 7 bits para selecionar o CHAR + 4 bits para escolher qual a LINHA dele
    output reg [7:0] data_font_rom  // saida: linha especifica do caractere especifico
);

reg [10:0] addr_reg;

always@(posedge dclk)
    addr_reg <= char_select;

always@*
    case (addr_reg)
        // code x00
        11'd0: data_font_rom = 8'b00000000; // 0
        11'd1: data_font_rom = 8'b00000000; // 1
        11'd2: data_font_rom = 8'b00000000; // 2
        11'd3: data_font_rom = 8'b00000000; // 3
        11'd4: data_font_rom = 8'b00000000; // 4
        11'd5: data_font_rom = 8'b00000000; // 5
        11'd6: data_font_rom = 8'b00000000; // 6
        11'd7: data_font_rom = 8'b00000000; // 7
        11'd8: data_font_rom = 8'b00000000; // 8
        11'd9: data_font_rom = 8'b00000000; // 9
        11'd10: data_font_rom = 8'b00000000; // a
        11'd11: data_font_rom = 8'b00000000; // b
        11'd12: data_font_rom = 8'b00000000; // c
        11'd13: data_font_rom = 8'b00000000; // d
        11'd14: data_font_rom = 8'b00000000; // e
        11'd15: data_font_rom = 8'b00000000; // f
        // code x01
        11'd16: data_font_rom = 8'b00000000; // 0
        11'd17: data_font_rom = 8'b00000000; // 1
        11'd18: data_font_rom = 8'b01111110; // 2  ******
        11'd19: data_font_rom = 8'b10000001; // 3 *      *
        11'd20: data_font_rom = 8'b10100101; // 4 * *  * *
        11'd21: data_font_rom = 8'b10000001; // 5 *      *
        11'd22: data_font_rom = 8'b10000001; // 6 *      *
        11'd23: data_font_rom = 8'b10111101; // 7 * **** *
        11'd24: data_font_rom = 8'b10011001; // 8 *  **  *
        11'd25: data_font_rom = 8'b10000001; // 9 *      *
        11'd26: data_font_rom = 8'b10000001; // a *      *
        11'd27: data_font_rom = 8'b01111110; // b  ******
        11'd28: data_font_rom = 8'b00000000; // c
        11'd29: data_font_rom = 8'b00000000; // d
        11'd30: data_font_rom = 8'b00000000; // e
        11'd31: data_font_rom = 8'b00000000; // f
        // code x02
        11'd32: data_font_rom = 8'b00000000; // 0
        11'd33: data_font_rom = 8'b00000000; // 1
        11'd34: data_font_rom = 8'b01111110; // 2  ******
        11'd35: data_font_rom = 8'b11111111; // 3 ********
        11'd36: data_font_rom = 8'b11011011; // 4 ** ** **
        11'd37: data_font_rom = 8'b11111111; // 5 ********
        11'd38: data_font_rom = 8'b11111111; // 6 ********
        11'd39: data_font_rom = 8'b11000011; // 7 **    **
        11'd40: data_font_rom = 8'b11100111; // 8 ***  ***
        11'd41: data_font_rom = 8'b11111111; // 9 ********
        11'd42: data_font_rom = 8'b11111111; // a ********
        11'd43: data_font_rom = 8'b01111110; // b  ******
        11'd44: data_font_rom = 8'b00000000; // c
        11'd45: data_font_rom = 8'b00000000; // d
        11'd46: data_font_rom = 8'b00000000; // e
        11'd47: data_font_rom = 8'b00000000; // f
        // code x03
        11'd48: data_font_rom = 8'b00000000; // 0
        11'd49: data_font_rom = 8'b00000000; // 1
        11'd50: data_font_rom = 8'b00000000; // 2
        11'd51: data_font_rom = 8'b00000000; // 3
        11'd52: data_font_rom = 8'b01101100; // 4  ** **
        11'd53: data_font_rom = 8'b11111110; // 5 *******
        11'd54: data_font_rom = 8'b11111110; // 6 *******
        11'd55: data_font_rom = 8'b11111110; // 7 *******
        11'd56: data_font_rom = 8'b11111110; // 8 *******
        11'd57: data_font_rom = 8'b01111100; // 9  *****
        11'd58: data_font_rom = 8'b00111000; // a   ***
        11'd59: data_font_rom = 8'b00010000; // b    *
        11'd60: data_font_rom = 8'b00000000; // c
        11'd61: data_font_rom = 8'b00000000; // d
        11'd62: data_font_rom = 8'b00000000; // e
        11'd63: data_font_rom = 8'b00000000; // f
        // code x04
        11'd64: data_font_rom = 8'b00000000; // 0
        11'd65: data_font_rom = 8'b00000000; // 1
        11'd66: data_font_rom = 8'b00000000; // 2
        11'd67: data_font_rom = 8'b00000000; // 3
        11'd68: data_font_rom = 8'b00010000; // 4    *
        11'd69: data_font_rom = 8'b00111000; // 5   ***
        11'd70: data_font_rom = 8'b01111100; // 6  *****
        11'd71: data_font_rom = 8'b11111110; // 7 *******
        11'd72: data_font_rom = 8'b01111100; // 8  *****
        11'd73: data_font_rom = 8'b00111000; // 9   ***
        11'd74: data_font_rom = 8'b00010000; // a    *
        11'd75: data_font_rom = 8'b00000000; // b
        11'd76: data_font_rom = 8'b00000000; // c
        11'd77: data_font_rom = 8'b00000000; // d
        11'd78: data_font_rom = 8'b00000000; // e
        11'd79: data_font_rom = 8'b00000000; // f
        // code x05
        11'd80: data_font_rom = 8'b00000000; // 0
        11'd81: data_font_rom = 8'b00000000; // 1
        11'd82: data_font_rom = 8'b00000000; // 2
        11'd83: data_font_rom = 8'b00011000; // 3    **
        11'd84: data_font_rom = 8'b00111100; // 4   ****
        11'd85: data_font_rom = 8'b00111100; // 5   ****
        11'd86: data_font_rom = 8'b11100111; // 6 ***  ***
        11'd87: data_font_rom = 8'b11100111; // 7 ***  ***
        11'd88: data_font_rom = 8'b11100111; // 8 ***  ***
        11'd89: data_font_rom = 8'b00011000; // 9    **
        11'd90: data_font_rom = 8'b00011000; // a    **
        11'd91: data_font_rom = 8'b00111100; // b   ****
        11'd92: data_font_rom = 8'b00000000; // c
        11'd93: data_font_rom = 8'b00000000; // d
        11'd94: data_font_rom = 8'b00000000; // e
        11'd95: data_font_rom = 8'b00000000; // f
        // code x06
        11'd96: data_font_rom = 8'b00000000; // 0
        11'd97: data_font_rom = 8'b00000000; // 1
        11'd98: data_font_rom = 8'b00000000; // 2
        11'd99: data_font_rom = 8'b00011000; // 3    **
        11'd100: data_font_rom = 8'b00111100; // 4   ****
        11'd101: data_font_rom = 8'b01111110; // 5  ******
        11'd102: data_font_rom = 8'b11111111; // 6 ********
        11'd103: data_font_rom = 8'b11111111; // 7 ********
        11'd104: data_font_rom = 8'b01111110; // 8  ******
        11'd105: data_font_rom = 8'b00011000; // 9    **
        11'd106: data_font_rom = 8'b00011000; // a    **
        11'd107: data_font_rom = 8'b00111100; // b   ****
        11'd108: data_font_rom = 8'b00000000; // c
        11'd109: data_font_rom = 8'b00000000; // d
        11'd110: data_font_rom = 8'b00000000; // e
        11'd111: data_font_rom = 8'b00000000; // f
        // code x07
        11'd112: data_font_rom = 8'b00000000; // 0
        11'd113: data_font_rom = 8'b00000000; // 1
        11'd114: data_font_rom = 8'b00000000; // 2
        11'd115: data_font_rom = 8'b00000000; // 3
        11'd116: data_font_rom = 8'b00000000; // 4
        11'd117: data_font_rom = 8'b00000000; // 5
        11'd118: data_font_rom = 8'b00011000; // 6    **
        11'd119: data_font_rom = 8'b00111100; // 7   ****
        11'd120: data_font_rom = 8'b00111100; // 8   ****
        11'd121: data_font_rom = 8'b00011000; // 9    **
        11'd122: data_font_rom = 8'b00000000; // a
        11'd123: data_font_rom = 8'b00000000; // b
        11'd124: data_font_rom = 8'b00000000; // c
        11'd125: data_font_rom = 8'b00000000; // d
        11'd126: data_font_rom = 8'b00000000; // e
        11'd127: data_font_rom = 8'b00000000; // f
        // code x08
        11'd128: data_font_rom = 8'b11111111; // 0 ********
        11'd129: data_font_rom = 8'b11111111; // 1 ********
        11'd130: data_font_rom = 8'b11111111; // 2 ********
        11'd131: data_font_rom = 8'b11111111; // 3 ********
        11'd132: data_font_rom = 8'b11111111; // 4 ********
        11'd133: data_font_rom = 8'b11111111; // 5 ********
        11'd134: data_font_rom = 8'b11100111; // 6 ***  ***
        11'd135: data_font_rom = 8'b11000011; // 7 **    **
        11'd136: data_font_rom = 8'b11000011; // 8 **    **
        11'd137: data_font_rom = 8'b11100111; // 9 ***  ***
        11'd138: data_font_rom = 8'b11111111; // a ********
        11'd139: data_font_rom = 8'b11111111; // b ********
        11'd140: data_font_rom = 8'b11111111; // c ********
        11'd141: data_font_rom = 8'b11111111; // d ********
        11'd142: data_font_rom = 8'b11111111; // e ********
        11'd143: data_font_rom = 8'b11111111; // f ********
        // code x09
        11'd144: data_font_rom = 8'b00000000; // 0
        11'd145: data_font_rom = 8'b00000000; // 1
        11'd146: data_font_rom = 8'b00000000; // 2
        11'd147: data_font_rom = 8'b00000000; // 3
        11'd148: data_font_rom = 8'b00000000; // 4
        11'd149: data_font_rom = 8'b00111100; // 5   ****
        11'd150: data_font_rom = 8'b01100110; // 6  **  **
        11'd151: data_font_rom = 8'b01000010; // 7  *    *
        11'd152: data_font_rom = 8'b01000010; // 8  *    *
        11'd153: data_font_rom = 8'b01100110; // 9  **  **
        11'd154: data_font_rom = 8'b00111100; // a   ****
        11'd155: data_font_rom = 8'b00000000; // b
        11'd156: data_font_rom = 8'b00000000; // c
        11'd157: data_font_rom = 8'b00000000; // d
        11'd158: data_font_rom = 8'b00000000; // e
        11'd159: data_font_rom = 8'b00000000; // f
        // code x0a
        11'd160: data_font_rom = 8'b11111111; // 0 ********
        11'd161: data_font_rom = 8'b11111111; // 1 ********
        11'd162: data_font_rom = 8'b11111111; // 2 ********
        11'd163: data_font_rom = 8'b11111111; // 3 ********
        11'd164: data_font_rom = 8'b11111111; // 4 ********
        11'd165: data_font_rom = 8'b11000011; // 5 **    **
        11'd166: data_font_rom = 8'b10011001; // 6 *  **  *
        11'd167: data_font_rom = 8'b10111101; // 7 * **** *
        11'd168: data_font_rom = 8'b10111101; // 8 * **** *
        11'd169: data_font_rom = 8'b10011001; // 9 *  **  *
        11'd170: data_font_rom = 8'b11000011; // a **    **
        11'd171: data_font_rom = 8'b11111111; // b ********
        11'd172: data_font_rom = 8'b11111111; // c ********
        11'd173: data_font_rom = 8'b11111111; // d ********
        11'd174: data_font_rom = 8'b11111111; // e ********
        11'd175: data_font_rom = 8'b11111111; // f ********
        // code x0b
        11'd176: data_font_rom = 8'b00000000; // 0
        11'd177: data_font_rom = 8'b00000000; // 1
        11'd178: data_font_rom = 8'b00011110; // 2    ****
        11'd179: data_font_rom = 8'b00001110; // 3     ***
        11'd180: data_font_rom = 8'b00011010; // 4    ** *
        11'd181: data_font_rom = 8'b00110010; // 5   **  *
        11'd182: data_font_rom = 8'b01111000; // 6  ****
        11'd183: data_font_rom = 8'b11001100; // 7 **  **
        11'd184: data_font_rom = 8'b11001100; // 8 **  **
        11'd185: data_font_rom = 8'b11001100; // 9 **  **
        11'd186: data_font_rom = 8'b11001100; // a **  **
        11'd187: data_font_rom = 8'b01111000; // b  ****
        11'd188: data_font_rom = 8'b00000000; // c
        11'd189: data_font_rom = 8'b00000000; // d
        11'd190: data_font_rom = 8'b00000000; // e
        11'd191: data_font_rom = 8'b00000000; // f
        // code x0c
        11'd192: data_font_rom = 8'b00000000; // 0
        11'd193: data_font_rom = 8'b00000000; // 1
        11'd194: data_font_rom = 8'b00111100; // 2   ****
        11'd195: data_font_rom = 8'b01100110; // 3  **  **
        11'd196: data_font_rom = 8'b01100110; // 4  **  **
        11'd197: data_font_rom = 8'b01100110; // 5  **  **
        11'd198: data_font_rom = 8'b01100110; // 6  **  **
        11'd199: data_font_rom = 8'b00111100; // 7   ****
        11'd200: data_font_rom = 8'b00011000; // 8    **
        11'd201: data_font_rom = 8'b01111110; // 9  ******
        11'd202: data_font_rom = 8'b00011000; // a    **
        11'd203: data_font_rom = 8'b00011000; // b    **
        11'd204: data_font_rom = 8'b00000000; // c
        11'd205: data_font_rom = 8'b00000000; // d
        11'd206: data_font_rom = 8'b00000000; // e
        11'd207: data_font_rom = 8'b00000000; // f
        // code x0d
        11'd208: data_font_rom = 8'b00000000; // 0
        11'd209: data_font_rom = 8'b00000000; // 1
        11'd210: data_font_rom = 8'b00111111; // 2   ******
        11'd211: data_font_rom = 8'b00110011; // 3   **  **
        11'd212: data_font_rom = 8'b00111111; // 4   ******
        11'd213: data_font_rom = 8'b00110000; // 5   **
        11'd214: data_font_rom = 8'b00110000; // 6   **
        11'd215: data_font_rom = 8'b00110000; // 7   **
        11'd216: data_font_rom = 8'b00110000; // 8   **
        11'd217: data_font_rom = 8'b01110000; // 9  ***
        11'd218: data_font_rom = 8'b11110000; // a ****
        11'd219: data_font_rom = 8'b11100000; // b ***
        11'd220: data_font_rom = 8'b00000000; // c
        11'd221: data_font_rom = 8'b00000000; // d
        11'd222: data_font_rom = 8'b00000000; // e
        11'd223: data_font_rom = 8'b00000000; // f
        // code x0e
        11'd224: data_font_rom = 8'b00000000; // 0
        11'd225: data_font_rom = 8'b00000000; // 1
        11'd226: data_font_rom = 8'b01111111; // 2  *******
        11'd227: data_font_rom = 8'b01100011; // 3  **   **
        11'd228: data_font_rom = 8'b01111111; // 4  *******
        11'd229: data_font_rom = 8'b01100011; // 5  **   **
        11'd230: data_font_rom = 8'b01100011; // 6  **   **
        11'd231: data_font_rom = 8'b01100011; // 7  **   **
        11'd232: data_font_rom = 8'b01100011; // 8  **   **
        11'd233: data_font_rom = 8'b01100111; // 9  **  ***
        11'd234: data_font_rom = 8'b11100111; // a ***  ***
        11'd235: data_font_rom = 8'b11100110; // b ***  **
        11'd236: data_font_rom = 8'b11000000; // c **
        11'd237: data_font_rom = 8'b00000000; // d
        11'd238: data_font_rom = 8'b00000000; // e
        11'd239: data_font_rom = 8'b00000000; // f
        // code x0f
        11'd240: data_font_rom = 8'b00000000; // 0
        11'd241: data_font_rom = 8'b00000000; // 1
        11'd242: data_font_rom = 8'b00000000; // 2
        11'd243: data_font_rom = 8'b00011000; // 3    **
        11'd244: data_font_rom = 8'b00011000; // 4    **
        11'd245: data_font_rom = 8'b11011011; // 5 ** ** **
        11'd246: data_font_rom = 8'b00111100; // 6   ****
        11'd247: data_font_rom = 8'b11100111; // 7 ***  ***
        11'd248: data_font_rom = 8'b00111100; // 8   ****
        11'd249: data_font_rom = 8'b11011011; // 9 ** ** **
        11'd250: data_font_rom = 8'b00011000; // a    **
        11'd251: data_font_rom = 8'b00011000; // b    **
        11'd252: data_font_rom = 8'b00000000; // c
        11'd253: data_font_rom = 8'b00000000; // d
        11'd254: data_font_rom = 8'b00000000; // e
        11'd255: data_font_rom = 8'b00000000; // f
        // code x10
        11'd256: data_font_rom = 8'b00000000; // 0
        11'd257: data_font_rom = 8'b10000000; // 1 *
        11'd258: data_font_rom = 8'b11000000; // 2 **
        11'd259: data_font_rom = 8'b11100000; // 3 ***
        11'd260: data_font_rom = 8'b11110000; // 4 ****
        11'd261: data_font_rom = 8'b11111000; // 5 *****
        11'd262: data_font_rom = 8'b11111110; // 6 *******
        11'd263: data_font_rom = 8'b11111000; // 7 *****
        11'd264: data_font_rom = 8'b11110000; // 8 ****
        11'd265: data_font_rom = 8'b11100000; // 9 ***
        11'd266: data_font_rom = 8'b11000000; // a **
        11'd267: data_font_rom = 8'b10000000; // b *
        11'd268: data_font_rom = 8'b00000000; // c
        11'd269: data_font_rom = 8'b00000000; // d
        11'd270: data_font_rom = 8'b00000000; // e
        11'd271: data_font_rom = 8'b00000000; // f
        // code x11
        11'd272: data_font_rom = 8'b00000000; // 0
        11'd273: data_font_rom = 8'b00000010; // 1       *
        11'd274: data_font_rom = 8'b00000110; // 2      **
        11'd275: data_font_rom = 8'b00001110; // 3     ***
        11'd276: data_font_rom = 8'b00011110; // 4    ****
        11'd277: data_font_rom = 8'b00111110; // 5   *****
        11'd278: data_font_rom = 8'b11111110; // 6 *******
        11'd279: data_font_rom = 8'b00111110; // 7   *****
        11'd280: data_font_rom = 8'b00011110; // 8    ****
        11'd281: data_font_rom = 8'b00001110; // 9     ***
        11'd282: data_font_rom = 8'b00000110; // a      **
        11'd283: data_font_rom = 8'b00000010; // b       *
        11'd284: data_font_rom = 8'b00000000; // c
        11'd285: data_font_rom = 8'b00000000; // d
        11'd286: data_font_rom = 8'b00000000; // e
        11'd287: data_font_rom = 8'b00000000; // f
        // code x12
        11'd288: data_font_rom = 8'b00000000; // 0
        11'd289: data_font_rom = 8'b00000000; // 1
        11'd290: data_font_rom = 8'b00011000; // 2    **
        11'd291: data_font_rom = 8'b00111100; // 3   ****
        11'd292: data_font_rom = 8'b01111110; // 4  ******
        11'd293: data_font_rom = 8'b00011000; // 5    **
        11'd294: data_font_rom = 8'b00011000; // 6    **
        11'd295: data_font_rom = 8'b00011000; // 7    **
        11'd296: data_font_rom = 8'b01111110; // 8  ******
        11'd297: data_font_rom = 8'b00111100; // 9   ****
        11'd298: data_font_rom = 8'b00011000; // a    **
        11'd299: data_font_rom = 8'b00000000; // b
        11'd300: data_font_rom = 8'b00000000; // c
        11'd301: data_font_rom = 8'b00000000; // d
        11'd302: data_font_rom = 8'b00000000; // e
        11'd303: data_font_rom = 8'b00000000; // f
        // code x13
        11'd304: data_font_rom = 8'b00000000; // 0
        11'd305: data_font_rom = 8'b00000000; // 1
        11'd306: data_font_rom = 8'b01100110; // 2  **  **
        11'd307: data_font_rom = 8'b01100110; // 3  **  **
        11'd308: data_font_rom = 8'b01100110; // 4  **  **
        11'd309: data_font_rom = 8'b01100110; // 5  **  **
        11'd310: data_font_rom = 8'b01100110; // 6  **  **
        11'd311: data_font_rom = 8'b01100110; // 7  **  **
        11'd312: data_font_rom = 8'b01100110; // 8  **  **
        11'd313: data_font_rom = 8'b00000000; // 9
        11'd314: data_font_rom = 8'b01100110; // a  **  **
        11'd315: data_font_rom = 8'b01100110; // b  **  **
        11'd316: data_font_rom = 8'b00000000; // c
        11'd317: data_font_rom = 8'b00000000; // d
        11'd318: data_font_rom = 8'b00000000; // e
        11'd319: data_font_rom = 8'b00000000; // f
        // code x14
        11'd320: data_font_rom = 8'b00000000; // 0
        11'd321: data_font_rom = 8'b00000000; // 1
        11'd322: data_font_rom = 8'b01111111; // 2  *******
        11'd323: data_font_rom = 8'b11011011; // 3 ** ** **
        11'd324: data_font_rom = 8'b11011011; // 4 ** ** **
        11'd325: data_font_rom = 8'b11011011; // 5 ** ** **
        11'd326: data_font_rom = 8'b01111011; // 6  **** **
        11'd327: data_font_rom = 8'b00011011; // 7    ** **
        11'd328: data_font_rom = 8'b00011011; // 8    ** **
        11'd329: data_font_rom = 8'b00011011; // 9    ** **
        11'd330: data_font_rom = 8'b00011011; // a    ** **
        11'd331: data_font_rom = 8'b00011011; // b    ** **
        11'd332: data_font_rom = 8'b00000000; // c
        11'd333: data_font_rom = 8'b00000000; // d
        11'd334: data_font_rom = 8'b00000000; // e
        11'd335: data_font_rom = 8'b00000000; // f
        // code x15
        11'd336: data_font_rom = 8'b00000000; // 0
        11'd337: data_font_rom = 8'b01111100; // 1  *****
        11'd338: data_font_rom = 8'b11000110; // 2 **   **
        11'd339: data_font_rom = 8'b01100000; // 3  **
        11'd340: data_font_rom = 8'b00111000; // 4   ***
        11'd341: data_font_rom = 8'b01101100; // 5  ** **
        11'd342: data_font_rom = 8'b11000110; // 6 **   **
        11'd343: data_font_rom = 8'b11000110; // 7 **   **
        11'd344: data_font_rom = 8'b01101100; // 8  ** **
        11'd345: data_font_rom = 8'b00111000; // 9   ***
        11'd346: data_font_rom = 8'b00001100; // a     **
        11'd347: data_font_rom = 8'b11000110; // b **   **
        11'd348: data_font_rom = 8'b01111100; // c  *****
        11'd349: data_font_rom = 8'b00000000; // d
        11'd350: data_font_rom = 8'b00000000; // e
        11'd351: data_font_rom = 8'b00000000; // f
        // code x16
        11'd352: data_font_rom = 8'b00000000; // 0
        11'd353: data_font_rom = 8'b00000000; // 1
        11'd354: data_font_rom = 8'b00000000; // 2
        11'd355: data_font_rom = 8'b00000000; // 3
        11'd356: data_font_rom = 8'b00000000; // 4
        11'd357: data_font_rom = 8'b00000000; // 5
        11'd358: data_font_rom = 8'b00000000; // 6
        11'd359: data_font_rom = 8'b00000000; // 7
        11'd360: data_font_rom = 8'b11111110; // 8 *******
        11'd361: data_font_rom = 8'b11111110; // 9 *******
        11'd362: data_font_rom = 8'b11111110; // a *******
        11'd363: data_font_rom = 8'b11111110; // b *******
        11'd364: data_font_rom = 8'b00000000; // c
        11'd365: data_font_rom = 8'b00000000; // d
        11'd366: data_font_rom = 8'b00000000; // e
        11'd367: data_font_rom = 8'b00000000; // f
        // code x17
        11'd368: data_font_rom = 8'b00000000; // 0
        11'd369: data_font_rom = 8'b00000000; // 1
        11'd370: data_font_rom = 8'b00011000; // 2    **
        11'd371: data_font_rom = 8'b00111100; // 3   ****
        11'd372: data_font_rom = 8'b01111110; // 4  ******
        11'd373: data_font_rom = 8'b00011000; // 5    **
        11'd374: data_font_rom = 8'b00011000; // 6    **
        11'd375: data_font_rom = 8'b00011000; // 7    **
        11'd376: data_font_rom = 8'b01111110; // 8  ******
        11'd377: data_font_rom = 8'b00111100; // 9   ****
        11'd378: data_font_rom = 8'b00011000; // a    **
        11'd379: data_font_rom = 8'b01111110; // b  ******
        11'd380: data_font_rom = 8'b00110000; // c
        11'd381: data_font_rom = 8'b00000000; // d
        11'd382: data_font_rom = 8'b00000000; // e
        11'd383: data_font_rom = 8'b00000000; // f
        // code x18
        11'd384: data_font_rom = 8'b00000000; // 0
        11'd385: data_font_rom = 8'b00000000; // 1
        11'd386: data_font_rom = 8'b00011000; // 2    **
        11'd387: data_font_rom = 8'b00111100; // 3   ****
        11'd388: data_font_rom = 8'b01111110; // 4  ******
        11'd389: data_font_rom = 8'b00011000; // 5    **
        11'd390: data_font_rom = 8'b00011000; // 6    **
        11'd391: data_font_rom = 8'b00011000; // 7    **
        11'd392: data_font_rom = 8'b00011000; // 8    **
        11'd393: data_font_rom = 8'b00011000; // 9    **
        11'd394: data_font_rom = 8'b00011000; // a    **
        11'd395: data_font_rom = 8'b00011000; // b    **
        11'd396: data_font_rom = 8'b00000000; // c
        11'd397: data_font_rom = 8'b00000000; // d
        11'd398: data_font_rom = 8'b00000000; // e
        11'd399: data_font_rom = 8'b00000000; // f
        // code x19
        11'd400: data_font_rom = 8'b00000000; // 0
        11'd401: data_font_rom = 8'b00000000; // 1
        11'd402: data_font_rom = 8'b00011000; // 2    **
        11'd403: data_font_rom = 8'b00011000; // 3    **
        11'd404: data_font_rom = 8'b00011000; // 4    **
        11'd405: data_font_rom = 8'b00011000; // 5    **
        11'd406: data_font_rom = 8'b00011000; // 6    **
        11'd407: data_font_rom = 8'b00011000; // 7    **
        11'd408: data_font_rom = 8'b00011000; // 8    **
        11'd409: data_font_rom = 8'b01111110; // 9  ******
        11'd410: data_font_rom = 8'b00111100; // a   ****
        11'd411: data_font_rom = 8'b00011000; // b    **
        11'd412: data_font_rom = 8'b00000000; // c
        11'd413: data_font_rom = 8'b00000000; // d
        11'd414: data_font_rom = 8'b00000000; // e
        11'd415: data_font_rom = 8'b00000000; // f
        // code x1a
        11'd416: data_font_rom = 8'b00000000; // 0
        11'd417: data_font_rom = 8'b00000000; // 1
        11'd418: data_font_rom = 8'b00000000; // 2
        11'd419: data_font_rom = 8'b00000000; // 3
        11'd420: data_font_rom = 8'b00000000; // 4
        11'd421: data_font_rom = 8'b00011000; // 5    **
        11'd422: data_font_rom = 8'b00001100; // 6     **
        11'd423: data_font_rom = 8'b11111110; // 7 *******
        11'd424: data_font_rom = 8'b00001100; // 8     **
        11'd425: data_font_rom = 8'b00011000; // 9    **
        11'd426: data_font_rom = 8'b00000000; // a
        11'd427: data_font_rom = 8'b00000000; // b
        11'd428: data_font_rom = 8'b00000000; // c
        11'd429: data_font_rom = 8'b00000000; // d
        11'd430: data_font_rom = 8'b00000000; // e
        11'd431: data_font_rom = 8'b00000000; // f
        // code x1b
        11'd432: data_font_rom = 8'b00000000; // 0
        11'd433: data_font_rom = 8'b00000000; // 1
        11'd434: data_font_rom = 8'b00000000; // 2
        11'd435: data_font_rom = 8'b00000000; // 3
        11'd436: data_font_rom = 8'b00000000; // 4
        11'd437: data_font_rom = 8'b00110000; // 5   **
        11'd438: data_font_rom = 8'b01100000; // 6  **
        11'd439: data_font_rom = 8'b11111110; // 7 *******
        11'd440: data_font_rom = 8'b01100000; // 8  **
        11'd441: data_font_rom = 8'b00110000; // 9   **
        11'd442: data_font_rom = 8'b00000000; // a
        11'd443: data_font_rom = 8'b00000000; // b
        11'd444: data_font_rom = 8'b00000000; // c
        11'd445: data_font_rom = 8'b00000000; // d
        11'd446: data_font_rom = 8'b00000000; // e
        11'd447: data_font_rom = 8'b00000000; // f
        // code x1c
        11'd448: data_font_rom = 8'b00000000; // 0
        11'd449: data_font_rom = 8'b00000000; // 1
        11'd450: data_font_rom = 8'b00000000; // 2
        11'd451: data_font_rom = 8'b00000000; // 3
        11'd452: data_font_rom = 8'b00000000; // 4
        11'd453: data_font_rom = 8'b00000000; // 5
        11'd454: data_font_rom = 8'b11000000; // 6 **
        11'd455: data_font_rom = 8'b11000000; // 7 **
        11'd456: data_font_rom = 8'b11000000; // 8 **
        11'd457: data_font_rom = 8'b11111110; // 9 *******
        11'd458: data_font_rom = 8'b00000000; // a
        11'd459: data_font_rom = 8'b00000000; // b
        11'd460: data_font_rom = 8'b00000000; // c
        11'd461: data_font_rom = 8'b00000000; // d
        11'd462: data_font_rom = 8'b00000000; // e
        11'd463: data_font_rom = 8'b00000000; // f
        // code x1d
        11'd464: data_font_rom = 8'b00000000; // 0
        11'd465: data_font_rom = 8'b00000000; // 1
        11'd466: data_font_rom = 8'b00000000; // 2
        11'd467: data_font_rom = 8'b00000000; // 3
        11'd468: data_font_rom = 8'b00000000; // 4
        11'd469: data_font_rom = 8'b00100100; // 5   *  *
        11'd470: data_font_rom = 8'b01100110; // 6  **  **
        11'd471: data_font_rom = 8'b11111111; // 7 ********
        11'd472: data_font_rom = 8'b01100110; // 8  **  **
        11'd473: data_font_rom = 8'b00100100; // 9   *  *
        11'd474: data_font_rom = 8'b00000000; // a
        11'd475: data_font_rom = 8'b00000000; // b
        11'd476: data_font_rom = 8'b00000000; // c
        11'd477: data_font_rom = 8'b00000000; // d
        11'd478: data_font_rom = 8'b00000000; // e
        11'd479: data_font_rom = 8'b00000000; // f
        // code x1e
        11'd480: data_font_rom = 8'b00000000; // 0
        11'd481: data_font_rom = 8'b00000000; // 1
        11'd482: data_font_rom = 8'b00000000; // 2
        11'd483: data_font_rom = 8'b00000000; // 3
        11'd484: data_font_rom = 8'b00010000; // 4    *
        11'd485: data_font_rom = 8'b00111000; // 5   ***
        11'd486: data_font_rom = 8'b00111000; // 6   ***
        11'd487: data_font_rom = 8'b01111100; // 7  *****
        11'd488: data_font_rom = 8'b01111100; // 8  *****
        11'd489: data_font_rom = 8'b11111110; // 9 *******
        11'd490: data_font_rom = 8'b11111110; // a *******
        11'd491: data_font_rom = 8'b00000000; // b
        11'd492: data_font_rom = 8'b00000000; // c
        11'd493: data_font_rom = 8'b00000000; // d
        11'd494: data_font_rom = 8'b00000000; // e
        11'd495: data_font_rom = 8'b00000000; // f
        // code x1f
        11'd496: data_font_rom = 8'b00000000; // 0
        11'd497: data_font_rom = 8'b00000000; // 1
        11'd498: data_font_rom = 8'b00000000; // 2
        11'd499: data_font_rom = 8'b00000000; // 3
        11'd500: data_font_rom = 8'b11111110; // 4 *******
        11'd501: data_font_rom = 8'b11111110; // 5 *******
        11'd502: data_font_rom = 8'b01111100; // 6  *****
        11'd503: data_font_rom = 8'b01111100; // 7  *****
        11'd504: data_font_rom = 8'b00111000; // 8   ***
        11'd505: data_font_rom = 8'b00111000; // 9   ***
        11'd506: data_font_rom = 8'b00010000; // a    *
        11'd507: data_font_rom = 8'b00000000; // b
        11'd508: data_font_rom = 8'b00000000; // c
        11'd509: data_font_rom = 8'b00000000; // d
        11'd510: data_font_rom = 8'b00000000; // e
        11'd511: data_font_rom = 8'b00000000; // f
        // code x20
        11'd512: data_font_rom = 8'b00000000; // 0
        11'd513: data_font_rom = 8'b00000000; // 1
        11'd514: data_font_rom = 8'b00000000; // 2
        11'd515: data_font_rom = 8'b00000000; // 3
        11'd516: data_font_rom = 8'b00000000; // 4
        11'd517: data_font_rom = 8'b00000000; // 5
        11'd518: data_font_rom = 8'b00000000; // 6
        11'd519: data_font_rom = 8'b00000000; // 7
        11'd520: data_font_rom = 8'b00000000; // 8
        11'd521: data_font_rom = 8'b00000000; // 9
        11'd522: data_font_rom = 8'b00000000; // a
        11'd523: data_font_rom = 8'b00000000; // b
        11'd524: data_font_rom = 8'b00000000; // c
        11'd525: data_font_rom = 8'b00000000; // d
        11'd526: data_font_rom = 8'b00000000; // e
        11'd527: data_font_rom = 8'b00000000; // f
        // code x21
        11'd528: data_font_rom = 8'b00000000; // 0
        11'd529: data_font_rom = 8'b00000000; // 1
        11'd530: data_font_rom = 8'b00011000; // 2    **
        11'd531: data_font_rom = 8'b00111100; // 3   ****
        11'd532: data_font_rom = 8'b00111100; // 4   ****
        11'd533: data_font_rom = 8'b00111100; // 5   ****
        11'd534: data_font_rom = 8'b00011000; // 6    **
        11'd535: data_font_rom = 8'b00011000; // 7    **
        11'd536: data_font_rom = 8'b00011000; // 8    **
        11'd537: data_font_rom = 8'b00000000; // 9
        11'd538: data_font_rom = 8'b00011000; // a    **
        11'd539: data_font_rom = 8'b00011000; // b    **
        11'd540: data_font_rom = 8'b00000000; // c
        11'd541: data_font_rom = 8'b00000000; // d
        11'd542: data_font_rom = 8'b00000000; // e
        11'd543: data_font_rom = 8'b00000000; // f
        // code x22
        11'd544: data_font_rom = 8'b00000000; // 0
        11'd545: data_font_rom = 8'b01100110; // 1  **  **
        11'd546: data_font_rom = 8'b01100110; // 2  **  **
        11'd547: data_font_rom = 8'b01100110; // 3  **  **
        11'd548: data_font_rom = 8'b00100100; // 4   *  *
        11'd549: data_font_rom = 8'b00000000; // 5
        11'd550: data_font_rom = 8'b00000000; // 6
        11'd551: data_font_rom = 8'b00000000; // 7
        11'd552: data_font_rom = 8'b00000000; // 8
        11'd553: data_font_rom = 8'b00000000; // 9
        11'd554: data_font_rom = 8'b00000000; // a
        11'd555: data_font_rom = 8'b00000000; // b
        11'd556: data_font_rom = 8'b00000000; // c
        11'd557: data_font_rom = 8'b00000000; // d
        11'd558: data_font_rom = 8'b00000000; // e
        11'd559: data_font_rom = 8'b00000000; // f
        // code x23
        11'd560: data_font_rom = 8'b00000000; // 0
        11'd561: data_font_rom = 8'b00000000; // 1
        11'd562: data_font_rom = 8'b00000000; // 2
        11'd563: data_font_rom = 8'b01101100; // 3  ** **
        11'd564: data_font_rom = 8'b01101100; // 4  ** **
        11'd565: data_font_rom = 8'b11111110; // 5 *******
        11'd566: data_font_rom = 8'b01101100; // 6  ** **
        11'd567: data_font_rom = 8'b01101100; // 7  ** **
        11'd568: data_font_rom = 8'b01101100; // 8  ** **
        11'd569: data_font_rom = 8'b11111110; // 9 *******
        11'd570: data_font_rom = 8'b01101100; // a  ** **
        11'd571: data_font_rom = 8'b01101100; // b  ** **
        11'd572: data_font_rom = 8'b00000000; // c
        11'd573: data_font_rom = 8'b00000000; // d
        11'd574: data_font_rom = 8'b00000000; // e
        11'd575: data_font_rom = 8'b00000000; // f
        // code x24
        11'd576: data_font_rom = 8'b00011000; // 0     **
        11'd577: data_font_rom = 8'b00011000; // 1     **
        11'd578: data_font_rom = 8'b01111100; // 2   *****
        11'd579: data_font_rom = 8'b11000110; // 3  **   **
        11'd580: data_font_rom = 8'b11000010; // 4  **    *
        11'd581: data_font_rom = 8'b11000000; // 5  **
        11'd582: data_font_rom = 8'b01111100; // 6   *****
        11'd583: data_font_rom = 8'b00000110; // 7       **
        11'd584: data_font_rom = 8'b00000110; // 8       **
        11'd585: data_font_rom = 8'b10000110; // 9  *    **
        11'd586: data_font_rom = 8'b11000110; // a  **   **
        11'd587: data_font_rom = 8'b01111100; // b   *****
        11'd588: data_font_rom = 8'b00011000; // c     **
        11'd589: data_font_rom = 8'b00011000; // d     **
        11'd590: data_font_rom = 8'b00000000; // e
        11'd591: data_font_rom = 8'b00000000; // f
        // code x25
        11'd592: data_font_rom = 8'b00000000; // 0
        11'd593: data_font_rom = 8'b00000000; // 1
        11'd594: data_font_rom = 8'b00000000; // 2
        11'd595: data_font_rom = 8'b00000000; // 3
        11'd596: data_font_rom = 8'b11000010; // 4 **    *
        11'd597: data_font_rom = 8'b11000110; // 5 **   **
        11'd598: data_font_rom = 8'b00001100; // 6     **
        11'd599: data_font_rom = 8'b00011000; // 7    **
        11'd600: data_font_rom = 8'b00110000; // 8   **
        11'd601: data_font_rom = 8'b01100000; // 9  **
        11'd602: data_font_rom = 8'b11000110; // a **   **
        11'd603: data_font_rom = 8'b10000110; // b *    **
        11'd604: data_font_rom = 8'b00000000; // c
        11'd605: data_font_rom = 8'b00000000; // d
        11'd606: data_font_rom = 8'b00000000; // e
        11'd607: data_font_rom = 8'b00000000; // f
        // code x26
        11'd608: data_font_rom = 8'b00000000; // 0
        11'd609: data_font_rom = 8'b00000000; // 1
        11'd610: data_font_rom = 8'b00111000; // 2   ***
        11'd611: data_font_rom = 8'b01101100; // 3  ** **
        11'd612: data_font_rom = 8'b01101100; // 4  ** **
        11'd613: data_font_rom = 8'b00111000; // 5   ***
        11'd614: data_font_rom = 8'b01110110; // 6  *** **
        11'd615: data_font_rom = 8'b11011100; // 7 ** ***
        11'd616: data_font_rom = 8'b11001100; // 8 **  **
        11'd617: data_font_rom = 8'b11001100; // 9 **  **
        11'd618: data_font_rom = 8'b11001100; // a **  **
        11'd619: data_font_rom = 8'b01110110; // b  *** **
        11'd620: data_font_rom = 8'b00000000; // c
        11'd621: data_font_rom = 8'b00000000; // d
        11'd622: data_font_rom = 8'b00000000; // e
        11'd623: data_font_rom = 8'b00000000; // f
        // code x27
        11'd624: data_font_rom = 8'b00000000; // 0
        11'd625: data_font_rom = 8'b00110000; // 1   **
        11'd626: data_font_rom = 8'b00110000; // 2   **
        11'd627: data_font_rom = 8'b00110000; // 3   **
        11'd628: data_font_rom = 8'b01100000; // 4  **
        11'd629: data_font_rom = 8'b00000000; // 5
        11'd630: data_font_rom = 8'b00000000; // 6
        11'd631: data_font_rom = 8'b00000000; // 7
        11'd632: data_font_rom = 8'b00000000; // 8
        11'd633: data_font_rom = 8'b00000000; // 9
        11'd634: data_font_rom = 8'b00000000; // a
        11'd635: data_font_rom = 8'b00000000; // b
        11'd636: data_font_rom = 8'b00000000; // c
        11'd637: data_font_rom = 8'b00000000; // d
        11'd638: data_font_rom = 8'b00000000; // e
        11'd639: data_font_rom = 8'b00000000; // f
        // code x28
        11'd640: data_font_rom = 8'b00000000; // 0
        11'd641: data_font_rom = 8'b00000000; // 1
        11'd642: data_font_rom = 8'b00001100; // 2     **
        11'd643: data_font_rom = 8'b00011000; // 3    **
        11'd644: data_font_rom = 8'b00110000; // 4   **
        11'd645: data_font_rom = 8'b00110000; // 5   **
        11'd646: data_font_rom = 8'b00110000; // 6   **
        11'd647: data_font_rom = 8'b00110000; // 7   **
        11'd648: data_font_rom = 8'b00110000; // 8   **
        11'd649: data_font_rom = 8'b00110000; // 9   **
        11'd650: data_font_rom = 8'b00011000; // a    **
        11'd651: data_font_rom = 8'b00001100; // b     **
        11'd652: data_font_rom = 8'b00000000; // c
        11'd653: data_font_rom = 8'b00000000; // d
        11'd654: data_font_rom = 8'b00000000; // e
        11'd655: data_font_rom = 8'b00000000; // f
        // code x29
        11'd656: data_font_rom = 8'b00000000; // 0
        11'd657: data_font_rom = 8'b00000000; // 1
        11'd658: data_font_rom = 8'b00110000; // 2   **
        11'd659: data_font_rom = 8'b00011000; // 3    **
        11'd660: data_font_rom = 8'b00001100; // 4     **
        11'd661: data_font_rom = 8'b00001100; // 5     **
        11'd662: data_font_rom = 8'b00001100; // 6     **
        11'd663: data_font_rom = 8'b00001100; // 7     **
        11'd664: data_font_rom = 8'b00001100; // 8     **
        11'd665: data_font_rom = 8'b00001100; // 9     **
        11'd666: data_font_rom = 8'b00011000; // a    **
        11'd667: data_font_rom = 8'b00110000; // b   **
        11'd668: data_font_rom = 8'b00000000; // c
        11'd669: data_font_rom = 8'b00000000; // d
        11'd670: data_font_rom = 8'b00000000; // e
        11'd671: data_font_rom = 8'b00000000; // f
        // code x2a
        11'd672: data_font_rom = 8'b00000000; // 0
        11'd673: data_font_rom = 8'b00000000; // 1
        11'd674: data_font_rom = 8'b00000000; // 2
        11'd675: data_font_rom = 8'b00000000; // 3
        11'd676: data_font_rom = 8'b00000000; // 4
        11'd677: data_font_rom = 8'b01100110; // 5  **  **
        11'd678: data_font_rom = 8'b00111100; // 6   ****
        11'd679: data_font_rom = 8'b11111111; // 7 ********
        11'd680: data_font_rom = 8'b00111100; // 8   ****
        11'd681: data_font_rom = 8'b01100110; // 9  **  **
        11'd682: data_font_rom = 8'b00000000; // a
        11'd683: data_font_rom = 8'b00000000; // b
        11'd684: data_font_rom = 8'b00000000; // c
        11'd685: data_font_rom = 8'b00000000; // d
        11'd686: data_font_rom = 8'b00000000; // e
        11'd687: data_font_rom = 8'b00000000; // f
        // code x2b
        11'd688: data_font_rom = 8'b00000000; // 0
        11'd689: data_font_rom = 8'b00000000; // 1
        11'd690: data_font_rom = 8'b00000000; // 2
        11'd691: data_font_rom = 8'b00000000; // 3
        11'd692: data_font_rom = 8'b00000000; // 4
        11'd693: data_font_rom = 8'b00011000; // 5    **
        11'd694: data_font_rom = 8'b00011000; // 6    **
        11'd695: data_font_rom = 8'b01111110; // 7  ******
        11'd696: data_font_rom = 8'b00011000; // 8    **
        11'd697: data_font_rom = 8'b00011000; // 9    **
        11'd698: data_font_rom = 8'b00000000; // a
        11'd699: data_font_rom = 8'b00000000; // b
        11'd700: data_font_rom = 8'b00000000; // c
        11'd701: data_font_rom = 8'b00000000; // d
        11'd702: data_font_rom = 8'b00000000; // e
        11'd703: data_font_rom = 8'b00000000; // f
        // code x2c
        11'd704: data_font_rom = 8'b00000000; // 0
        11'd705: data_font_rom = 8'b00000000; // 1
        11'd706: data_font_rom = 8'b00000000; // 2
        11'd707: data_font_rom = 8'b00000000; // 3
        11'd708: data_font_rom = 8'b00000000; // 4
        11'd709: data_font_rom = 8'b00000000; // 5
        11'd710: data_font_rom = 8'b00000000; // 6
        11'd711: data_font_rom = 8'b00000000; // 7
        11'd712: data_font_rom = 8'b00000000; // 8
        11'd713: data_font_rom = 8'b00011000; // 9    **
        11'd714: data_font_rom = 8'b00011000; // a    **
        11'd715: data_font_rom = 8'b00011000; // b    **
        11'd716: data_font_rom = 8'b00110000; // c   **
        11'd717: data_font_rom = 8'b00000000; // d
        11'd718: data_font_rom = 8'b00000000; // e
        11'd719: data_font_rom = 8'b00000000; // f
        // code x2d
        11'd720: data_font_rom = 8'b00000000; // 0
        11'd721: data_font_rom = 8'b00000000; // 1
        11'd722: data_font_rom = 8'b00000000; // 2
        11'd723: data_font_rom = 8'b00000000; // 3
        11'd724: data_font_rom = 8'b00000000; // 4
        11'd725: data_font_rom = 8'b00000000; // 5
        11'd726: data_font_rom = 8'b00000000; // 6
        11'd727: data_font_rom = 8'b01111110; // 7  ******
        11'd728: data_font_rom = 8'b00000000; // 8
        11'd729: data_font_rom = 8'b00000000; // 9
        11'd730: data_font_rom = 8'b00000000; // a
        11'd731: data_font_rom = 8'b00000000; // b
        11'd732: data_font_rom = 8'b00000000; // c
        11'd733: data_font_rom = 8'b00000000; // d
        11'd734: data_font_rom = 8'b00000000; // e
        11'd735: data_font_rom = 8'b00000000; // f
        // code x2e
        11'd736: data_font_rom = 8'b00000000; // 0
        11'd737: data_font_rom = 8'b00000000; // 1
        11'd738: data_font_rom = 8'b00000000; // 2
        11'd739: data_font_rom = 8'b00000000; // 3
        11'd740: data_font_rom = 8'b00000000; // 4
        11'd741: data_font_rom = 8'b00000000; // 5
        11'd742: data_font_rom = 8'b00000000; // 6
        11'd743: data_font_rom = 8'b00000000; // 7
        11'd744: data_font_rom = 8'b00000000; // 8
        11'd745: data_font_rom = 8'b00000000; // 9
        11'd746: data_font_rom = 8'b00011000; // a    **
        11'd747: data_font_rom = 8'b00011000; // b    **
        11'd748: data_font_rom = 8'b00000000; // c
        11'd749: data_font_rom = 8'b00000000; // d
        11'd750: data_font_rom = 8'b00000000; // e
        11'd751: data_font_rom = 8'b00000000; // f
        // code x2f
        11'd752: data_font_rom = 8'b00000000; // 0
        11'd753: data_font_rom = 8'b00000000; // 1
        11'd754: data_font_rom = 8'b00000000; // 2
        11'd755: data_font_rom = 8'b00000000; // 3
        11'd756: data_font_rom = 8'b00000010; // 4       *
        11'd757: data_font_rom = 8'b00000110; // 5      **
        11'd758: data_font_rom = 8'b00001100; // 6     **
        11'd759: data_font_rom = 8'b00011000; // 7    **
        11'd760: data_font_rom = 8'b00110000; // 8   **
        11'd761: data_font_rom = 8'b01100000; // 9  **
        11'd762: data_font_rom = 8'b11000000; // a **
        11'd763: data_font_rom = 8'b10000000; // b *
        11'd764: data_font_rom = 8'b00000000; // c
        11'd765: data_font_rom = 8'b00000000; // d
        11'd766: data_font_rom = 8'b00000000; // e
        11'd767: data_font_rom = 8'b00000000; // f
        // code x30
        11'd768: data_font_rom = 8'b00000000; // 0
        11'd769: data_font_rom = 8'b00000000; // 1
        11'd770: data_font_rom = 8'b01111100; // 2  *****
        11'd771: data_font_rom = 8'b11000110; // 3 **   **
        11'd772: data_font_rom = 8'b11000110; // 4 **   **
        11'd773: data_font_rom = 8'b11001110; // 5 **  ***
        11'd774: data_font_rom = 8'b11011110; // 6 ** ****
        11'd775: data_font_rom = 8'b11110110; // 7 **** **
        11'd776: data_font_rom = 8'b11100110; // 8 ***  **
        11'd777: data_font_rom = 8'b11000110; // 9 **   **
        11'd778: data_font_rom = 8'b11000110; // a **   **
        11'd779: data_font_rom = 8'b01111100; // b  *****
        11'd780: data_font_rom = 8'b00000000; // c
        11'd781: data_font_rom = 8'b00000000; // d
        11'd782: data_font_rom = 8'b00000000; // e
        11'd783: data_font_rom = 8'b00000000; // f
        // code x31
        11'd784: data_font_rom = 8'b00000000; // 0
        11'd785: data_font_rom = 8'b00000000; // 1
        11'd786: data_font_rom = 8'b00011000; // 2
        11'd787: data_font_rom = 8'b00111000; // 3
        11'd788: data_font_rom = 8'b01111000; // 4    **
        11'd789: data_font_rom = 8'b00011000; // 5   ***
        11'd790: data_font_rom = 8'b00011000; // 6  ****
        11'd791: data_font_rom = 8'b00011000; // 7    **
        11'd792: data_font_rom = 8'b00011000; // 8    **
        11'd793: data_font_rom = 8'b00011000; // 9    **
        11'd794: data_font_rom = 8'b00011000; // a    **
        11'd795: data_font_rom = 8'b01111110; // b    **
        11'd796: data_font_rom = 8'b00000000; // c    **
        11'd797: data_font_rom = 8'b00000000; // d  ******
        11'd798: data_font_rom = 8'b00000000; // e
        11'd799: data_font_rom = 8'b00000000; // f
        // code x32
        11'd800: data_font_rom = 8'b00000000; // 0
        11'd801: data_font_rom = 8'b00000000; // 1
        11'd802: data_font_rom = 8'b01111100; // 2  *****
        11'd803: data_font_rom = 8'b11000110; // 3 **   **
        11'd804: data_font_rom = 8'b00000110; // 4      **
        11'd805: data_font_rom = 8'b00001100; // 5     **
        11'd806: data_font_rom = 8'b00011000; // 6    **
        11'd807: data_font_rom = 8'b00110000; // 7   **
        11'd808: data_font_rom = 8'b01100000; // 8  **
        11'd809: data_font_rom = 8'b11000000; // 9 **
        11'd810: data_font_rom = 8'b11000110; // a **   **
        11'd811: data_font_rom = 8'b11111110; // b *******
        11'd812: data_font_rom = 8'b00000000; // c
        11'd813: data_font_rom = 8'b00000000; // d
        11'd814: data_font_rom = 8'b00000000; // e
        11'd815: data_font_rom = 8'b00000000; // f
        // code x33
        11'd816: data_font_rom = 8'b00000000; // 0
        11'd817: data_font_rom = 8'b00000000; // 1
        11'd818: data_font_rom = 8'b01111100; // 2  *****
        11'd819: data_font_rom = 8'b11000110; // 3 **   **
        11'd820: data_font_rom = 8'b00000110; // 4      **
        11'd821: data_font_rom = 8'b00000110; // 5      **
        11'd822: data_font_rom = 8'b00111100; // 6   ****
        11'd823: data_font_rom = 8'b00000110; // 7      **
        11'd824: data_font_rom = 8'b00000110; // 8      **
        11'd825: data_font_rom = 8'b00000110; // 9      **
        11'd826: data_font_rom = 8'b11000110; // a **   **
        11'd827: data_font_rom = 8'b01111100; // b  *****
        11'd828: data_font_rom = 8'b00000000; // c
        11'd829: data_font_rom = 8'b00000000; // d
        11'd830: data_font_rom = 8'b00000000; // e
        11'd831: data_font_rom = 8'b00000000; // f
        // code x34
        11'd832: data_font_rom = 8'b00000000; // 0
        11'd833: data_font_rom = 8'b00000000; // 1
        11'd834: data_font_rom = 8'b00001100; // 2     **
        11'd835: data_font_rom = 8'b00011100; // 3    ***
        11'd836: data_font_rom = 8'b00111100; // 4   ****
        11'd837: data_font_rom = 8'b01101100; // 5  ** **
        11'd838: data_font_rom = 8'b11001100; // 6 **  **
        11'd839: data_font_rom = 8'b11111110; // 7 *******
        11'd840: data_font_rom = 8'b00001100; // 8     **
        11'd841: data_font_rom = 8'b00001100; // 9     **
        11'd842: data_font_rom = 8'b00001100; // a     **
        11'd843: data_font_rom = 8'b00011110; // b    ****
        11'd844: data_font_rom = 8'b00000000; // c
        11'd845: data_font_rom = 8'b00000000; // d
        11'd846: data_font_rom = 8'b00000000; // e
        11'd847: data_font_rom = 8'b00000000; // f
        // code x35
        11'd848: data_font_rom = 8'b00000000; // 0
        11'd849: data_font_rom = 8'b00000000; // 1
        11'd850: data_font_rom = 8'b11111110; // 2 *******
        11'd851: data_font_rom = 8'b11000000; // 3 **
        11'd852: data_font_rom = 8'b11000000; // 4 **
        11'd853: data_font_rom = 8'b11000000; // 5 **
        11'd854: data_font_rom = 8'b11111100; // 6 ******
        11'd855: data_font_rom = 8'b00000110; // 7      **
        11'd856: data_font_rom = 8'b00000110; // 8      **
        11'd857: data_font_rom = 8'b00000110; // 9      **
        11'd858: data_font_rom = 8'b11000110; // a **   **
        11'd859: data_font_rom = 8'b01111100; // b  *****
        11'd860: data_font_rom = 8'b00000000; // c
        11'd861: data_font_rom = 8'b00000000; // d
        11'd862: data_font_rom = 8'b00000000; // e
        11'd863: data_font_rom = 8'b00000000; // f
        // code x36
        11'd864: data_font_rom = 8'b00000000; // 0
        11'd865: data_font_rom = 8'b00000000; // 1
        11'd866: data_font_rom = 8'b00111000; // 2   ***
        11'd867: data_font_rom = 8'b01100000; // 3  **
        11'd868: data_font_rom = 8'b11000000; // 4 **
        11'd869: data_font_rom = 8'b11000000; // 5 **
        11'd870: data_font_rom = 8'b11111100; // 6 ******
        11'd871: data_font_rom = 8'b11000110; // 7 **   **
        11'd872: data_font_rom = 8'b11000110; // 8 **   **
        11'd873: data_font_rom = 8'b11000110; // 9 **   **
        11'd874: data_font_rom = 8'b11000110; // a **   **
        11'd875: data_font_rom = 8'b01111100; // b  *****
        11'd876: data_font_rom = 8'b00000000; // c
        11'd877: data_font_rom = 8'b00000000; // d
        11'd878: data_font_rom = 8'b00000000; // e
        11'd879: data_font_rom = 8'b00000000; // f
        // code x37
        11'd880: data_font_rom = 8'b00000000; // 0
        11'd881: data_font_rom = 8'b00000000; // 1
        11'd882: data_font_rom = 8'b11111110; // 2 *******
        11'd883: data_font_rom = 8'b11000110; // 3 **   **
        11'd884: data_font_rom = 8'b00000110; // 4      **
        11'd885: data_font_rom = 8'b00000110; // 5      **
        11'd886: data_font_rom = 8'b00001100; // 6     **
        11'd887: data_font_rom = 8'b00011000; // 7    **
        11'd888: data_font_rom = 8'b00110000; // 8   **
        11'd889: data_font_rom = 8'b00110000; // 9   **
        11'd890: data_font_rom = 8'b00110000; // a   **
        11'd891: data_font_rom = 8'b00110000; // b   **
        11'd892: data_font_rom = 8'b00000000; // c
        11'd893: data_font_rom = 8'b00000000; // d
        11'd894: data_font_rom = 8'b00000000; // e
        11'd895: data_font_rom = 8'b00000000; // f
        // code x38
        11'd896: data_font_rom = 8'b00000000; // 0
        11'd897: data_font_rom = 8'b00000000; // 1
        11'd898: data_font_rom = 8'b01111100; // 2  *****
        11'd899: data_font_rom = 8'b11000110; // 3 **   **
        11'd900: data_font_rom = 8'b11000110; // 4 **   **
        11'd901: data_font_rom = 8'b11000110; // 5 **   **
        11'd902: data_font_rom = 8'b01111100; // 6  *****
        11'd903: data_font_rom = 8'b11000110; // 7 **   **
        11'd904: data_font_rom = 8'b11000110; // 8 **   **
        11'd905: data_font_rom = 8'b11000110; // 9 **   **
        11'd906: data_font_rom = 8'b11000110; // a **   **
        11'd907: data_font_rom = 8'b01111100; // b  *****
        11'd908: data_font_rom = 8'b00000000; // c
        11'd909: data_font_rom = 8'b00000000; // d
        11'd910: data_font_rom = 8'b00000000; // e
        11'd911: data_font_rom = 8'b00000000; // f
        // code x39
        11'd912: data_font_rom = 8'b00000000; // 0
        11'd913: data_font_rom = 8'b00000000; // 1
        11'd914: data_font_rom = 8'b01111100; // 2  *****
        11'd915: data_font_rom = 8'b11000110; // 3 **   **
        11'd916: data_font_rom = 8'b11000110; // 4 **   **
        11'd917: data_font_rom = 8'b11000110; // 5 **   **
        11'd918: data_font_rom = 8'b01111110; // 6  ******
        11'd919: data_font_rom = 8'b00000110; // 7      **
        11'd920: data_font_rom = 8'b00000110; // 8      **
        11'd921: data_font_rom = 8'b00000110; // 9      **
        11'd922: data_font_rom = 8'b00001100; // a     **
        11'd923: data_font_rom = 8'b01111000; // b  ****
        11'd924: data_font_rom = 8'b00000000; // c
        11'd925: data_font_rom = 8'b00000000; // d
        11'd926: data_font_rom = 8'b00000000; // e
        11'd927: data_font_rom = 8'b00000000; // f
        // code x3a
        11'd928: data_font_rom = 8'b00000000; // 0
        11'd929: data_font_rom = 8'b00000000; // 1
        11'd930: data_font_rom = 8'b00000000; // 2
        11'd931: data_font_rom = 8'b00000000; // 3
        11'd932: data_font_rom = 8'b00011000; // 4    **
        11'd933: data_font_rom = 8'b00011000; // 5    **
        11'd934: data_font_rom = 8'b00000000; // 6
        11'd935: data_font_rom = 8'b00000000; // 7
        11'd936: data_font_rom = 8'b00000000; // 8
        11'd937: data_font_rom = 8'b00011000; // 9    **
        11'd938: data_font_rom = 8'b00011000; // a    **
        11'd939: data_font_rom = 8'b00000000; // b
        11'd940: data_font_rom = 8'b00000000; // c
        11'd941: data_font_rom = 8'b00000000; // d
        11'd942: data_font_rom = 8'b00000000; // e
        11'd943: data_font_rom = 8'b00000000; // f
        // code x3b
        11'd944: data_font_rom = 8'b00000000; // 0
        11'd945: data_font_rom = 8'b00000000; // 1
        11'd946: data_font_rom = 8'b00000000; // 2
        11'd947: data_font_rom = 8'b00000000; // 3
        11'd948: data_font_rom = 8'b00011000; // 4    **
        11'd949: data_font_rom = 8'b00011000; // 5    **
        11'd950: data_font_rom = 8'b00000000; // 6
        11'd951: data_font_rom = 8'b00000000; // 7
        11'd952: data_font_rom = 8'b00000000; // 8
        11'd953: data_font_rom = 8'b00011000; // 9    **
        11'd954: data_font_rom = 8'b00011000; // a    **
        11'd955: data_font_rom = 8'b00110000; // b   **
        11'd956: data_font_rom = 8'b00000000; // c
        11'd957: data_font_rom = 8'b00000000; // d
        11'd958: data_font_rom = 8'b00000000; // e
        11'd959: data_font_rom = 8'b00000000; // f
        // code x3c
        11'd960: data_font_rom = 8'b00000000; // 0
        11'd961: data_font_rom = 8'b00000000; // 1
        11'd962: data_font_rom = 8'b00000000; // 2
        11'd963: data_font_rom = 8'b00000110; // 3      **
        11'd964: data_font_rom = 8'b00001100; // 4     **
        11'd965: data_font_rom = 8'b00011000; // 5    **
        11'd966: data_font_rom = 8'b00110000; // 6   **
        11'd967: data_font_rom = 8'b01100000; // 7  **
        11'd968: data_font_rom = 8'b00110000; // 8   **
        11'd969: data_font_rom = 8'b00011000; // 9    **
        11'd970: data_font_rom = 8'b00001100; // a     **
        11'd971: data_font_rom = 8'b00000110; // b      **
        11'd972: data_font_rom = 8'b00000000; // c
        11'd973: data_font_rom = 8'b00000000; // d
        11'd974: data_font_rom = 8'b00000000; // e
        11'd975: data_font_rom = 8'b00000000; // f
        // code x3d
        11'd976: data_font_rom = 8'b00000000; // 0
        11'd977: data_font_rom = 8'b00000000; // 1
        11'd978: data_font_rom = 8'b00000000; // 2
        11'd979: data_font_rom = 8'b00000000; // 3
        11'd980: data_font_rom = 8'b00000000; // 4
        11'd981: data_font_rom = 8'b01111110; // 5  ******
        11'd982: data_font_rom = 8'b00000000; // 6
        11'd983: data_font_rom = 8'b00000000; // 7
        11'd984: data_font_rom = 8'b01111110; // 8  ******
        11'd985: data_font_rom = 8'b00000000; // 9
        11'd986: data_font_rom = 8'b00000000; // a
        11'd987: data_font_rom = 8'b00000000; // b
        11'd988: data_font_rom = 8'b00000000; // c
        11'd989: data_font_rom = 8'b00000000; // d
        11'd990: data_font_rom = 8'b00000000; // e
        11'd991: data_font_rom = 8'b00000000; // f
        // code x3e
        11'd992: data_font_rom = 8'b00000000; // 0
        11'd993: data_font_rom = 8'b00000000; // 1
        11'd994: data_font_rom = 8'b00000000; // 2
        11'd995: data_font_rom = 8'b01100000; // 3  **
        11'd996: data_font_rom = 8'b00110000; // 4   **
        11'd997: data_font_rom = 8'b00011000; // 5    **
        11'd998: data_font_rom = 8'b00001100; // 6     **
        11'd999: data_font_rom = 8'b00000110; // 7      **
        11'd1000: data_font_rom = 8'b00001100; // 8     **
        11'd1001: data_font_rom = 8'b00011000; // 9    **
        11'd1002: data_font_rom = 8'b00110000; // a   **
        11'd1003: data_font_rom = 8'b01100000; // b  **
        11'd1004: data_font_rom = 8'b00000000; // c
        11'd1005: data_font_rom = 8'b00000000; // d
        11'd1006: data_font_rom = 8'b00000000; // e
        11'd1007: data_font_rom = 8'b00000000; // f
        // code x3f
        11'd1008: data_font_rom = 8'b00000000; // 0
        11'd1009: data_font_rom = 8'b00000000; // 1
        11'd1010: data_font_rom = 8'b01111100; // 2  *****
        11'd1011: data_font_rom = 8'b11000110; // 3 **   **
        11'd1012: data_font_rom = 8'b11000110; // 4 **   **
        11'd1013: data_font_rom = 8'b00001100; // 5     **
        11'd1014: data_font_rom = 8'b00011000; // 6    **
        11'd1015: data_font_rom = 8'b00011000; // 7    **
        11'd1016: data_font_rom = 8'b00011000; // 8    **
        11'd1017: data_font_rom = 8'b00000000; // 9
        11'd1018: data_font_rom = 8'b00011000; // a    **
        11'd1019: data_font_rom = 8'b00011000; // b    **
        11'd1020: data_font_rom = 8'b00000000; // c
        11'd1021: data_font_rom = 8'b00000000; // d
        11'd1022: data_font_rom = 8'b00000000; // e
        11'd1023: data_font_rom = 8'b00000000; // f
        // code x40
        11'd1024: data_font_rom = 8'b00000000; // 0
        11'd1025: data_font_rom = 8'b00000000; // 1
        11'd1026: data_font_rom = 8'b01111100; // 2  *****
        11'd1027: data_font_rom = 8'b11000110; // 3 **   **
        11'd1028: data_font_rom = 8'b11000110; // 4 **   **
        11'd1029: data_font_rom = 8'b11000110; // 5 **   **
        11'd1030: data_font_rom = 8'b11011110; // 6 ** ****
        11'd1031: data_font_rom = 8'b11011110; // 7 ** ****
        11'd1032: data_font_rom = 8'b11011110; // 8 ** ****
        11'd1033: data_font_rom = 8'b11011100; // 9 ** ***
        11'd1034: data_font_rom = 8'b11000000; // a **
        11'd1035: data_font_rom = 8'b01111100; // b  *****
        11'd1036: data_font_rom = 8'b00000000; // c
        11'd1037: data_font_rom = 8'b00000000; // d
        11'd1038: data_font_rom = 8'b00000000; // e
        11'd1039: data_font_rom = 8'b00000000; // f
        // code x41
        11'd1040: data_font_rom = 8'b00000000; // 0
        11'd1041: data_font_rom = 8'b00000000; // 1
        11'd1042: data_font_rom = 8'b00010000; // 2    *
        11'd1043: data_font_rom = 8'b00111000; // 3   ***
        11'd1044: data_font_rom = 8'b01101100; // 4  ** **
        11'd1045: data_font_rom = 8'b11000110; // 5 **   **
        11'd1046: data_font_rom = 8'b11000110; // 6 **   **
        11'd1047: data_font_rom = 8'b11111110; // 7 *******
        11'd1048: data_font_rom = 8'b11000110; // 8 **   **
        11'd1049: data_font_rom = 8'b11000110; // 9 **   **
        11'd1050: data_font_rom = 8'b11000110; // a **   **
        11'd1051: data_font_rom = 8'b11000110; // b **   **
        11'd1052: data_font_rom = 8'b00000000; // c
        11'd1053: data_font_rom = 8'b00000000; // d
        11'd1054: data_font_rom = 8'b00000000; // e
        11'd1055: data_font_rom = 8'b00000000; // f
        // code x42
        11'd1056: data_font_rom = 8'b00000000; // 0
        11'd1057: data_font_rom = 8'b00000000; // 1
        11'd1058: data_font_rom = 8'b11111100; // 2 ******
        11'd1059: data_font_rom = 8'b01100110; // 3  **  **
        11'd1060: data_font_rom = 8'b01100110; // 4  **  **
        11'd1061: data_font_rom = 8'b01100110; // 5  **  **
        11'd1062: data_font_rom = 8'b01111100; // 6  *****
        11'd1063: data_font_rom = 8'b01100110; // 7  **  **
        11'd1064: data_font_rom = 8'b01100110; // 8  **  **
        11'd1065: data_font_rom = 8'b01100110; // 9  **  **
        11'd1066: data_font_rom = 8'b01100110; // a  **  **
        11'd1067: data_font_rom = 8'b11111100; // b ******
        11'd1068: data_font_rom = 8'b00000000; // c
        11'd1069: data_font_rom = 8'b00000000; // d
        11'd1070: data_font_rom = 8'b00000000; // e
        11'd1071: data_font_rom = 8'b00000000; // f
        // code x43
        11'd1072: data_font_rom = 8'b00000000; // 0
        11'd1073: data_font_rom = 8'b00000000; // 1
        11'd1074: data_font_rom = 8'b00111100; // 2   ****
        11'd1075: data_font_rom = 8'b01100110; // 3  **  **
        11'd1076: data_font_rom = 8'b11000010; // 4 **    *
        11'd1077: data_font_rom = 8'b11000000; // 5 **
        11'd1078: data_font_rom = 8'b11000000; // 6 **
        11'd1079: data_font_rom = 8'b11000000; // 7 **
        11'd1080: data_font_rom = 8'b11000000; // 8 **
        11'd1081: data_font_rom = 8'b11000010; // 9 **    *
        11'd1082: data_font_rom = 8'b01100110; // a  **  **
        11'd1083: data_font_rom = 8'b00111100; // b   ****
        11'd1084: data_font_rom = 8'b00000000; // c
        11'd1085: data_font_rom = 8'b00000000; // d
        11'd1086: data_font_rom = 8'b00000000; // e
        11'd1087: data_font_rom = 8'b00000000; // f
        // code x44
        11'd1088: data_font_rom = 8'b00000000; // 0
        11'd1089: data_font_rom = 8'b00000000; // 1
        11'd1090: data_font_rom = 8'b11111000; // 2 *****
        11'd1091: data_font_rom = 8'b01101100; // 3  ** **
        11'd1092: data_font_rom = 8'b01100110; // 4  **  **
        11'd1093: data_font_rom = 8'b01100110; // 5  **  **
        11'd1094: data_font_rom = 8'b01100110; // 6  **  **
        11'd1095: data_font_rom = 8'b01100110; // 7  **  **
        11'd1096: data_font_rom = 8'b01100110; // 8  **  **
        11'd1097: data_font_rom = 8'b01100110; // 9  **  **
        11'd1098: data_font_rom = 8'b01101100; // a  ** **
        11'd1099: data_font_rom = 8'b11111000; // b *****
        11'd1100: data_font_rom = 8'b00000000; // c
        11'd1101: data_font_rom = 8'b00000000; // d
        11'd1102: data_font_rom = 8'b00000000; // e
        11'd1103: data_font_rom = 8'b00000000; // f
        // code x45
        11'd1104: data_font_rom = 8'b00000000; // 0
        11'd1105: data_font_rom = 8'b00000000; // 1
        11'd1106: data_font_rom = 8'b11111110; // 2 *******
        11'd1107: data_font_rom = 8'b01100110; // 3  **  **
        11'd1108: data_font_rom = 8'b01100010; // 4  **   *
        11'd1109: data_font_rom = 8'b01101000; // 5  ** *
        11'd1110: data_font_rom = 8'b01111000; // 6  ****
        11'd1111: data_font_rom = 8'b01101000; // 7  ** *
        11'd1112: data_font_rom = 8'b01100000; // 8  **
        11'd1113: data_font_rom = 8'b01100010; // 9  **   *
        11'd1114: data_font_rom = 8'b01100110; // a  **  **
        11'd1115: data_font_rom = 8'b11111110; // b *******
        11'd1116: data_font_rom = 8'b00000000; // c
        11'd1117: data_font_rom = 8'b00000000; // d
        11'd1118: data_font_rom = 8'b00000000; // e
        11'd1119: data_font_rom = 8'b00000000; // f
        // code x46
        11'd1120: data_font_rom = 8'b00000000; // 0
        11'd1121: data_font_rom = 8'b00000000; // 1
        11'd1122: data_font_rom = 8'b11111110; // 2 *******
        11'd1123: data_font_rom = 8'b01100110; // 3  **  **
        11'd1124: data_font_rom = 8'b01100010; // 4  **   *
        11'd1125: data_font_rom = 8'b01101000; // 5  ** *
        11'd1126: data_font_rom = 8'b01111000; // 6  ****
        11'd1127: data_font_rom = 8'b01101000; // 7  ** *
        11'd1128: data_font_rom = 8'b01100000; // 8  **
        11'd1129: data_font_rom = 8'b01100000; // 9  **
        11'd1130: data_font_rom = 8'b01100000; // a  **
        11'd1131: data_font_rom = 8'b11110000; // b ****
        11'd1132: data_font_rom = 8'b00000000; // c
        11'd1133: data_font_rom = 8'b00000000; // d
        11'd1134: data_font_rom = 8'b00000000; // e
        11'd1135: data_font_rom = 8'b00000000; // f
        // code x47
        11'd1136: data_font_rom = 8'b00000000; // 0
        11'd1137: data_font_rom = 8'b00000000; // 1
        11'd1138: data_font_rom = 8'b00111100; // 2   ****
        11'd1139: data_font_rom = 8'b01100110; // 3  **  **
        11'd1140: data_font_rom = 8'b11000010; // 4 **    *
        11'd1141: data_font_rom = 8'b11000000; // 5 **
        11'd1142: data_font_rom = 8'b11000000; // 6 **
        11'd1143: data_font_rom = 8'b11011110; // 7 ** ****
        11'd1144: data_font_rom = 8'b11000110; // 8 **   **
        11'd1145: data_font_rom = 8'b11000110; // 9 **   **
        11'd1146: data_font_rom = 8'b01100110; // a  **  **
        11'd1147: data_font_rom = 8'b00111010; // b   *** *
        11'd1148: data_font_rom = 8'b00000000; // c
        11'd1149: data_font_rom = 8'b00000000; // d
        11'd1150: data_font_rom = 8'b00000000; // e
        11'd1151: data_font_rom = 8'b00000000; // f
        // code x48
        11'd1152: data_font_rom = 8'b00000000; // 0
        11'd1153: data_font_rom = 8'b00000000; // 1
        11'd1154: data_font_rom = 8'b11000110; // 2 **   **
        11'd1155: data_font_rom = 8'b11000110; // 3 **   **
        11'd1156: data_font_rom = 8'b11000110; // 4 **   **
        11'd1157: data_font_rom = 8'b11000110; // 5 **   **
        11'd1158: data_font_rom = 8'b11111110; // 6 *******
        11'd1159: data_font_rom = 8'b11000110; // 7 **   **
        11'd1160: data_font_rom = 8'b11000110; // 8 **   **
        11'd1161: data_font_rom = 8'b11000110; // 9 **   **
        11'd1162: data_font_rom = 8'b11000110; // a **   **
        11'd1163: data_font_rom = 8'b11000110; // b **   **
        11'd1164: data_font_rom = 8'b00000000; // c
        11'd1165: data_font_rom = 8'b00000000; // d
        11'd1166: data_font_rom = 8'b00000000; // e
        11'd1167: data_font_rom = 8'b00000000; // f
        // code x49
        11'd1168: data_font_rom = 8'b00000000; // 0
        11'd1169: data_font_rom = 8'b00000000; // 1
        11'd1170: data_font_rom = 8'b00111100; // 2   ****
        11'd1171: data_font_rom = 8'b00011000; // 3    **
        11'd1172: data_font_rom = 8'b00011000; // 4    **
        11'd1173: data_font_rom = 8'b00011000; // 5    **
        11'd1174: data_font_rom = 8'b00011000; // 6    **
        11'd1175: data_font_rom = 8'b00011000; // 7    **
        11'd1176: data_font_rom = 8'b00011000; // 8    **
        11'd1177: data_font_rom = 8'b00011000; // 9    **
        11'd1178: data_font_rom = 8'b00011000; // a    **
        11'd1179: data_font_rom = 8'b00111100; // b   ****
        11'd1180: data_font_rom = 8'b00000000; // c
        11'd1181: data_font_rom = 8'b00000000; // d
        11'd1182: data_font_rom = 8'b00000000; // e
        11'd1183: data_font_rom = 8'b00000000; // f
        // code x4a
        11'd1184: data_font_rom = 8'b00000000; // 0
        11'd1185: data_font_rom = 8'b00000000; // 1
        11'd1186: data_font_rom = 8'b00011110; // 2    ****
        11'd1187: data_font_rom = 8'b00001100; // 3     **
        11'd1188: data_font_rom = 8'b00001100; // 4     **
        11'd1189: data_font_rom = 8'b00001100; // 5     **
        11'd1190: data_font_rom = 8'b00001100; // 6     **
        11'd1191: data_font_rom = 8'b00001100; // 7     **
        11'd1192: data_font_rom = 8'b11001100; // 8 **  **
        11'd1193: data_font_rom = 8'b11001100; // 9 **  **
        11'd1194: data_font_rom = 8'b11001100; // a **  **
        11'd1195: data_font_rom = 8'b01111000; // b  ****
        11'd1196: data_font_rom = 8'b00000000; // c
        11'd1197: data_font_rom = 8'b00000000; // d
        11'd1198: data_font_rom = 8'b00000000; // e
        11'd1199: data_font_rom = 8'b00000000; // f
        // code x4b
        11'd1200: data_font_rom = 8'b00000000; // 0
        11'd1201: data_font_rom = 8'b00000000; // 1
        11'd1202: data_font_rom = 8'b11100110; // 2 ***  **
        11'd1203: data_font_rom = 8'b01100110; // 3  **  **
        11'd1204: data_font_rom = 8'b01100110; // 4  **  **
        11'd1205: data_font_rom = 8'b01101100; // 5  ** **
        11'd1206: data_font_rom = 8'b01111000; // 6  ****
        11'd1207: data_font_rom = 8'b01111000; // 7  ****
        11'd1208: data_font_rom = 8'b01101100; // 8  ** **
        11'd1209: data_font_rom = 8'b01100110; // 9  **  **
        11'd1210: data_font_rom = 8'b01100110; // a  **  **
        11'd1211: data_font_rom = 8'b11100110; // b ***  **
        11'd1212: data_font_rom = 8'b00000000; // c
        11'd1213: data_font_rom = 8'b00000000; // d
        11'd1214: data_font_rom = 8'b00000000; // e
        11'd1215: data_font_rom = 8'b00000000; // f
        // code x4c
        11'd1216: data_font_rom = 8'b00000000; // 0
        11'd1217: data_font_rom = 8'b00000000; // 1
        11'd1218: data_font_rom = 8'b11110000; // 2 ****
        11'd1219: data_font_rom = 8'b01100000; // 3  **
        11'd1220: data_font_rom = 8'b01100000; // 4  **
        11'd1221: data_font_rom = 8'b01100000; // 5  **
        11'd1222: data_font_rom = 8'b01100000; // 6  **
        11'd1223: data_font_rom = 8'b01100000; // 7  **
        11'd1224: data_font_rom = 8'b01100000; // 8  **
        11'd1225: data_font_rom = 8'b01100010; // 9  **   *
        11'd1226: data_font_rom = 8'b01100110; // a  **  **
        11'd1227: data_font_rom = 8'b11111110; // b *******
        11'd1228: data_font_rom = 8'b00000000; // c
        11'd1229: data_font_rom = 8'b00000000; // d
        11'd1230: data_font_rom = 8'b00000000; // e
        11'd1231: data_font_rom = 8'b00000000; // f
        // code x4d
        11'd1232: data_font_rom = 8'b00000000; // 0
        11'd1233: data_font_rom = 8'b00000000; // 1
        11'd1234: data_font_rom = 8'b11000011; // 2 **    **
        11'd1235: data_font_rom = 8'b11100111; // 3 ***  ***
        11'd1236: data_font_rom = 8'b11111111; // 4 ********
        11'd1237: data_font_rom = 8'b11111111; // 5 ********
        11'd1238: data_font_rom = 8'b11011011; // 6 ** ** **
        11'd1239: data_font_rom = 8'b11000011; // 7 **    **
        11'd1240: data_font_rom = 8'b11000011; // 8 **    **
        11'd1241: data_font_rom = 8'b11000011; // 9 **    **
        11'd1242: data_font_rom = 8'b11000011; // a **    **
        11'd1243: data_font_rom = 8'b11000011; // b **    **
        11'd1244: data_font_rom = 8'b00000000; // c
        11'd1245: data_font_rom = 8'b00000000; // d
        11'd1246: data_font_rom = 8'b00000000; // e
        11'd1247: data_font_rom = 8'b00000000; // f
        // code x4e
        11'd1248: data_font_rom = 8'b00000000; // 0
        11'd1249: data_font_rom = 8'b00000000; // 1
        11'd1250: data_font_rom = 8'b11000110; // 2 **   **
        11'd1251: data_font_rom = 8'b11100110; // 3 ***  **
        11'd1252: data_font_rom = 8'b11110110; // 4 **** **
        11'd1253: data_font_rom = 8'b11111110; // 5 *******
        11'd1254: data_font_rom = 8'b11011110; // 6 ** ****
        11'd1255: data_font_rom = 8'b11001110; // 7 **  ***
        11'd1256: data_font_rom = 8'b11000110; // 8 **   **
        11'd1257: data_font_rom = 8'b11000110; // 9 **   **
        11'd1258: data_font_rom = 8'b11000110; // a **   **
        11'd1259: data_font_rom = 8'b11000110; // b **   **
        11'd1260: data_font_rom = 8'b00000000; // c
        11'd1261: data_font_rom = 8'b00000000; // d
        11'd1262: data_font_rom = 8'b00000000; // e
        11'd1263: data_font_rom = 8'b00000000; // f
        // code x4f
        11'd1264: data_font_rom = 8'b00000000; // 0
        11'd1265: data_font_rom = 8'b00000000; // 1
        11'd1266: data_font_rom = 8'b01111100; // 2  *****
        11'd1267: data_font_rom = 8'b11000110; // 3 **   **
        11'd1268: data_font_rom = 8'b11000110; // 4 **   **
        11'd1269: data_font_rom = 8'b11000110; // 5 **   **
        11'd1270: data_font_rom = 8'b11000110; // 6 **   **
        11'd1271: data_font_rom = 8'b11000110; // 7 **   **
        11'd1272: data_font_rom = 8'b11000110; // 8 **   **
        11'd1273: data_font_rom = 8'b11000110; // 9 **   **
        11'd1274: data_font_rom = 8'b11000110; // a **   **
        11'd1275: data_font_rom = 8'b01111100; // b  *****
        11'd1276: data_font_rom = 8'b00000000; // c
        11'd1277: data_font_rom = 8'b00000000; // d
        11'd1278: data_font_rom = 8'b00000000; // e
        11'd1279: data_font_rom = 8'b00000000; // f
        // code x50
        11'd1280: data_font_rom = 8'b00000000; // 0
        11'd1281: data_font_rom = 8'b00000000; // 1
        11'd1282: data_font_rom = 8'b11111100; // 2 ******
        11'd1283: data_font_rom = 8'b01100110; // 3  **  **
        11'd1284: data_font_rom = 8'b01100110; // 4  **  **
        11'd1285: data_font_rom = 8'b01100110; // 5  **  **
        11'd1286: data_font_rom = 8'b01111100; // 6  *****
        11'd1287: data_font_rom = 8'b01100000; // 7  **
        11'd1288: data_font_rom = 8'b01100000; // 8  **
        11'd1289: data_font_rom = 8'b01100000; // 9  **
        11'd1290: data_font_rom = 8'b01100000; // a  **
        11'd1291: data_font_rom = 8'b11110000; // b ****
        11'd1292: data_font_rom = 8'b00000000; // c
        11'd1293: data_font_rom = 8'b00000000; // d
        11'd1294: data_font_rom = 8'b00000000; // e
        11'd1295: data_font_rom = 8'b00000000; // f
        // code x510
        11'd1296: data_font_rom = 8'b00000000; // 0
        11'd1297: data_font_rom = 8'b00000000; // 1
        11'd1298: data_font_rom = 8'b01111100; // 2  *****
        11'd1299: data_font_rom = 8'b11000110; // 3 **   **
        11'd1300: data_font_rom = 8'b11000110; // 4 **   **
        11'd1301: data_font_rom = 8'b11000110; // 5 **   **
        11'd1302: data_font_rom = 8'b11000110; // 6 **   **
        11'd1303: data_font_rom = 8'b11000110; // 7 **   **
        11'd1304: data_font_rom = 8'b11000110; // 8 **   **
        11'd1305: data_font_rom = 8'b11010110; // 9 ** * **
        11'd1306: data_font_rom = 8'b11011110; // a ** ****
        11'd1307: data_font_rom = 8'b01111100; // b  *****
        11'd1308: data_font_rom = 8'b00001100; // c     **
        11'd1309: data_font_rom = 8'b00001110; // d     ***
        11'd1310: data_font_rom = 8'b00000000; // e
        11'd1311: data_font_rom = 8'b00000000; // f
        // code x52
        11'd1312: data_font_rom = 8'b00000000; // 0
        11'd1313: data_font_rom = 8'b00000000; // 1
        11'd1314: data_font_rom = 8'b11111100; // 2 ******
        11'd1315: data_font_rom = 8'b01100110; // 3  **  **
        11'd1316: data_font_rom = 8'b01100110; // 4  **  **
        11'd1317: data_font_rom = 8'b01100110; // 5  **  **
        11'd1318: data_font_rom = 8'b01111100; // 6  *****
        11'd1319: data_font_rom = 8'b01101100; // 7  ** **
        11'd1320: data_font_rom = 8'b01100110; // 8  **  **
        11'd1321: data_font_rom = 8'b01100110; // 9  **  **
        11'd1322: data_font_rom = 8'b01100110; // a  **  **
        11'd1323: data_font_rom = 8'b11100110; // b ***  **
        11'd1324: data_font_rom = 8'b00000000; // c
        11'd1325: data_font_rom = 8'b00000000; // d
        11'd1326: data_font_rom = 8'b00000000; // e
        11'd1327: data_font_rom = 8'b00000000; // f
        // code x53
        11'd1328: data_font_rom = 8'b00000000; // 0
        11'd1329: data_font_rom = 8'b00000000; // 1
        11'd1330: data_font_rom = 8'b01111100; // 2  *****
        11'd1331: data_font_rom = 8'b11000110; // 3 **   **
        11'd1332: data_font_rom = 8'b11000110; // 4 **   **
        11'd1333: data_font_rom = 8'b01100000; // 5  **
        11'd1334: data_font_rom = 8'b00111000; // 6   ***
        11'd1335: data_font_rom = 8'b00001100; // 7     **
        11'd1336: data_font_rom = 8'b00000110; // 8      **
        11'd1337: data_font_rom = 8'b11000110; // 9 **   **
        11'd1338: data_font_rom = 8'b11000110; // a **   **
        11'd1339: data_font_rom = 8'b01111100; // b  *****
        11'd1340: data_font_rom = 8'b00000000; // c
        11'd1341: data_font_rom = 8'b00000000; // d
        11'd1342: data_font_rom = 8'b00000000; // e
        11'd1343: data_font_rom = 8'b00000000; // f
        // code x54
        11'd1344: data_font_rom = 8'b00000000; // 0
        11'd1345: data_font_rom = 8'b00000000; // 1
        11'd1346: data_font_rom = 8'b11111111; // 2 ********
        11'd1347: data_font_rom = 8'b11011011; // 3 ** ** **
        11'd1348: data_font_rom = 8'b10011001; // 4 *  **  *
        11'd1349: data_font_rom = 8'b00011000; // 5    **
        11'd1350: data_font_rom = 8'b00011000; // 6    **
        11'd1351: data_font_rom = 8'b00011000; // 7    **
        11'd1352: data_font_rom = 8'b00011000; // 8    **
        11'd1353: data_font_rom = 8'b00011000; // 9    **
        11'd1354: data_font_rom = 8'b00011000; // a    **
        11'd1355: data_font_rom = 8'b00111100; // b   ****
        11'd1356: data_font_rom = 8'b00000000; // c
        11'd1357: data_font_rom = 8'b00000000; // d
        11'd1358: data_font_rom = 8'b00000000; // e
        11'd1359: data_font_rom = 8'b00000000; // f
        // code x55
        11'd1360: data_font_rom = 8'b00000000; // 0
        11'd1361: data_font_rom = 8'b00000000; // 1
        11'd1362: data_font_rom = 8'b11000110; // 2 **   **
        11'd1363: data_font_rom = 8'b11000110; // 3 **   **
        11'd1364: data_font_rom = 8'b11000110; // 4 **   **
        11'd1365: data_font_rom = 8'b11000110; // 5 **   **
        11'd1366: data_font_rom = 8'b11000110; // 6 **   **
        11'd1367: data_font_rom = 8'b11000110; // 7 **   **
        11'd1368: data_font_rom = 8'b11000110; // 8 **   **
        11'd1369: data_font_rom = 8'b11000110; // 9 **   **
        11'd1370: data_font_rom = 8'b11000110; // a **   **
        11'd1371: data_font_rom = 8'b01111100; // b  *****
        11'd1372: data_font_rom = 8'b00000000; // c
        11'd1373: data_font_rom = 8'b00000000; // d
        11'd1374: data_font_rom = 8'b00000000; // e
        11'd1375: data_font_rom = 8'b00000000; // f
        // code x56
        11'd1376: data_font_rom = 8'b00000000; // 0
        11'd1377: data_font_rom = 8'b00000000; // 1
        11'd1378: data_font_rom = 8'b11000011; // 2 **    **
        11'd1379: data_font_rom = 8'b11000011; // 3 **    **
        11'd1380: data_font_rom = 8'b11000011; // 4 **    **
        11'd1381: data_font_rom = 8'b11000011; // 5 **    **
        11'd1382: data_font_rom = 8'b11000011; // 6 **    **
        11'd1383: data_font_rom = 8'b11000011; // 7 **    **
        11'd1384: data_font_rom = 8'b11000011; // 8 **    **
        11'd1385: data_font_rom = 8'b01100110; // 9  **  **
        11'd1386: data_font_rom = 8'b00111100; // a   ****
        11'd1387: data_font_rom = 8'b00011000; // b    **
        11'd1388: data_font_rom = 8'b00000000; // c
        11'd1389: data_font_rom = 8'b00000000; // d
        11'd1390: data_font_rom = 8'b00000000; // e
        11'd1391: data_font_rom = 8'b00000000; // f
        // code x57
        11'd1392: data_font_rom = 8'b00000000; // 0
        11'd1393: data_font_rom = 8'b00000000; // 1
        11'd1394: data_font_rom = 8'b11000011; // 2 **    **
        11'd1395: data_font_rom = 8'b11000011; // 3 **    **
        11'd1396: data_font_rom = 8'b11000011; // 4 **    **
        11'd1397: data_font_rom = 8'b11000011; // 5 **    **
        11'd1398: data_font_rom = 8'b11000011; // 6 **    **
        11'd1399: data_font_rom = 8'b11011011; // 7 ** ** **
        11'd1400: data_font_rom = 8'b11011011; // 8 ** ** **
        11'd1401: data_font_rom = 8'b11111111; // 9 ********
        11'd1402: data_font_rom = 8'b01100110; // a  **  **
        11'd1403: data_font_rom = 8'b01100110; // b  **  **
        11'd1404: data_font_rom = 8'b00000000; // c
        11'd1405: data_font_rom = 8'b00000000; // d
        11'd1406: data_font_rom = 8'b00000000; // e
        11'd1407: data_font_rom = 8'b00000000; // f
        // code x58
        11'd1408: data_font_rom = 8'b00000000; // 0
        11'd1409: data_font_rom = 8'b00000000; // 1
        11'd1410: data_font_rom = 8'b11000011; // 2 **    **
        11'd1411: data_font_rom = 8'b11000011; // 3 **    **
        11'd1412: data_font_rom = 8'b01100110; // 4  **  **
        11'd1413: data_font_rom = 8'b00111100; // 5   ****
        11'd1414: data_font_rom = 8'b00011000; // 6    **
        11'd1415: data_font_rom = 8'b00011000; // 7    **
        11'd1416: data_font_rom = 8'b00111100; // 8   ****
        11'd1417: data_font_rom = 8'b01100110; // 9  **  **
        11'd1418: data_font_rom = 8'b11000011; // a **    **
        11'd1419: data_font_rom = 8'b11000011; // b **    **
        11'd1420: data_font_rom = 8'b00000000; // c
        11'd1421: data_font_rom = 8'b00000000; // d
        11'd1422: data_font_rom = 8'b00000000; // e
        11'd1423: data_font_rom = 8'b00000000; // f
        // code x59
        11'd1424: data_font_rom = 8'b00000000; // 0
        11'd1425: data_font_rom = 8'b00000000; // 1
        11'd1426: data_font_rom = 8'b11000011; // 2 **    **
        11'd1427: data_font_rom = 8'b11000011; // 3 **    **
        11'd1428: data_font_rom = 8'b11000011; // 4 **    **
        11'd1429: data_font_rom = 8'b01100110; // 5  **  **
        11'd1430: data_font_rom = 8'b00111100; // 6   ****
        11'd1431: data_font_rom = 8'b00011000; // 7    **
        11'd1432: data_font_rom = 8'b00011000; // 8    **
        11'd1433: data_font_rom = 8'b00011000; // 9    **
        11'd1434: data_font_rom = 8'b00011000; // a    **
        11'd1435: data_font_rom = 8'b00111100; // b   ****
        11'd1436: data_font_rom = 8'b00000000; // c
        11'd1437: data_font_rom = 8'b00000000; // d
        11'd1438: data_font_rom = 8'b00000000; // e
        11'd1439: data_font_rom = 8'b00000000; // f
        // code x5a
        11'd1440: data_font_rom = 8'b00000000; // 0
        11'd1441: data_font_rom = 8'b00000000; // 1
        11'd1442: data_font_rom = 8'b11111111; // 2 ********
        11'd1443: data_font_rom = 8'b11000011; // 3 **    **
        11'd1444: data_font_rom = 8'b10000110; // 4 *    **
        11'd1445: data_font_rom = 8'b00001100; // 5     **
        11'd1446: data_font_rom = 8'b00011000; // 6    **
        11'd1447: data_font_rom = 8'b00110000; // 7   **
        11'd1448: data_font_rom = 8'b01100000; // 8  **
        11'd1449: data_font_rom = 8'b11000001; // 9 **     *
        11'd1450: data_font_rom = 8'b11000011; // a **    **
        11'd1451: data_font_rom = 8'b11111111; // b ********
        11'd1452: data_font_rom = 8'b00000000; // c
        11'd1453: data_font_rom = 8'b00000000; // d
        11'd1454: data_font_rom = 8'b00000000; // e
        11'd1455: data_font_rom = 8'b00000000; // f
        // code x5b
        11'd1456: data_font_rom = 8'b00000000; // 0
        11'd1457: data_font_rom = 8'b00000000; // 1
        11'd1458: data_font_rom = 8'b00111100; // 2   ****
        11'd1459: data_font_rom = 8'b00110000; // 3   **
        11'd1460: data_font_rom = 8'b00110000; // 4   **
        11'd1461: data_font_rom = 8'b00110000; // 5   **
        11'd1462: data_font_rom = 8'b00110000; // 6   **
        11'd1463: data_font_rom = 8'b00110000; // 7   **
        11'd1464: data_font_rom = 8'b00110000; // 8   **
        11'd1465: data_font_rom = 8'b00110000; // 9   **
        11'd1466: data_font_rom = 8'b00110000; // a   **
        11'd1467: data_font_rom = 8'b00111100; // b   ****
        11'd1468: data_font_rom = 8'b00000000; // c
        11'd1469: data_font_rom = 8'b00000000; // d
        11'd1470: data_font_rom = 8'b00000000; // e
        11'd1471: data_font_rom = 8'b00000000; // f
        // code x5c
        11'd1472: data_font_rom = 8'b00000000; // 0
        11'd1473: data_font_rom = 8'b00000000; // 1
        11'd1474: data_font_rom = 8'b00000000; // 2
        11'd1475: data_font_rom = 8'b10000000; // 3 *
        11'd1476: data_font_rom = 8'b11000000; // 4 **
        11'd1477: data_font_rom = 8'b11100000; // 5 ***
        11'd1478: data_font_rom = 8'b01110000; // 6  ***
        11'd1479: data_font_rom = 8'b00111000; // 7   ***
        11'd1480: data_font_rom = 8'b00011100; // 8    ***
        11'd1481: data_font_rom = 8'b00001110; // 9     ***
        11'd1482: data_font_rom = 8'b00000110; // a      **
        11'd1483: data_font_rom = 8'b00000010; // b       *
        11'd1484: data_font_rom = 8'b00000000; // c
        11'd1485: data_font_rom = 8'b00000000; // d
        11'd1486: data_font_rom = 8'b00000000; // e
        11'd1487: data_font_rom = 8'b00000000; // f
        // code x5d
        11'd1488: data_font_rom = 8'b00000000; // 0
        11'd1489: data_font_rom = 8'b00000000; // 1
        11'd1490: data_font_rom = 8'b00111100; // 2   ****
        11'd1491: data_font_rom = 8'b00001100; // 3     **
        11'd1492: data_font_rom = 8'b00001100; // 4     **
        11'd1493: data_font_rom = 8'b00001100; // 5     **
        11'd1494: data_font_rom = 8'b00001100; // 6     **
        11'd1495: data_font_rom = 8'b00001100; // 7     **
        11'd1496: data_font_rom = 8'b00001100; // 8     **
        11'd1497: data_font_rom = 8'b00001100; // 9     **
        11'd1498: data_font_rom = 8'b00001100; // a     **
        11'd1499: data_font_rom = 8'b00111100; // b   ****
        11'd1500: data_font_rom = 8'b00000000; // c
        11'd1501: data_font_rom = 8'b00000000; // d
        11'd1502: data_font_rom = 8'b00000000; // e
        11'd1503: data_font_rom = 8'b00000000; // f
        // code x5e
        11'd1504: data_font_rom = 8'b00010000; // 0    *
        11'd1505: data_font_rom = 8'b00111000; // 1   ***
        11'd1506: data_font_rom = 8'b01101100; // 2  ** **
        11'd1507: data_font_rom = 8'b11000110; // 3 **   **
        11'd1508: data_font_rom = 8'b00000000; // 4
        11'd1509: data_font_rom = 8'b00000000; // 5
        11'd1510: data_font_rom = 8'b00000000; // 6
        11'd1511: data_font_rom = 8'b00000000; // 7
        11'd1512: data_font_rom = 8'b00000000; // 8
        11'd1513: data_font_rom = 8'b00000000; // 9
        11'd1514: data_font_rom = 8'b00000000; // a
        11'd1515: data_font_rom = 8'b00000000; // b
        11'd1516: data_font_rom = 8'b00000000; // c
        11'd1517: data_font_rom = 8'b00000000; // d
        11'd1518: data_font_rom = 8'b00000000; // e
        11'd1519: data_font_rom = 8'b00000000; // f
        // code x5f
        11'd1520: data_font_rom = 8'b00000000; // 0
        11'd1521: data_font_rom = 8'b00000000; // 1
        11'd1522: data_font_rom = 8'b00000000; // 2
        11'd1523: data_font_rom = 8'b00000000; // 3
        11'd1524: data_font_rom = 8'b00000000; // 4
        11'd1525: data_font_rom = 8'b00000000; // 5
        11'd1526: data_font_rom = 8'b00000000; // 6
        11'd1527: data_font_rom = 8'b00000000; // 7
        11'd1528: data_font_rom = 8'b00000000; // 8
        11'd1529: data_font_rom = 8'b00000000; // 9
        11'd1530: data_font_rom = 8'b00000000; // a
        11'd1531: data_font_rom = 8'b00000000; // b
        11'd1532: data_font_rom = 8'b00000000; // c
        11'd1533: data_font_rom = 8'b11111111; // d ********
        11'd1534: data_font_rom = 8'b00000000; // e
        11'd1535: data_font_rom = 8'b00000000; // f
        // code x60
        11'd1536: data_font_rom = 8'b00110000; // 0   **
        11'd1537: data_font_rom = 8'b00110000; // 1   **
        11'd1538: data_font_rom = 8'b00011000; // 2    **
        11'd1539: data_font_rom = 8'b00000000; // 3
        11'd1540: data_font_rom = 8'b00000000; // 4
        11'd1541: data_font_rom = 8'b00000000; // 5
        11'd1542: data_font_rom = 8'b00000000; // 6
        11'd1543: data_font_rom = 8'b00000000; // 7
        11'd1544: data_font_rom = 8'b00000000; // 8
        11'd1545: data_font_rom = 8'b00000000; // 9
        11'd1546: data_font_rom = 8'b00000000; // a
        11'd1547: data_font_rom = 8'b00000000; // b
        11'd1548: data_font_rom = 8'b00000000; // c
        11'd1549: data_font_rom = 8'b00000000; // d
        11'd1550: data_font_rom = 8'b00000000; // e
        11'd1551: data_font_rom = 8'b00000000; // f
        // code x61
        11'd1552: data_font_rom = 8'b00000000; // 0
        11'd1553: data_font_rom = 8'b00000000; // 1
        11'd1554: data_font_rom = 8'b00000000; // 2
        11'd1555: data_font_rom = 8'b00000000; // 3
        11'd1556: data_font_rom = 8'b00000000; // 4
        11'd1557: data_font_rom = 8'b01111000; // 5  ****
        11'd1558: data_font_rom = 8'b00001100; // 6     **
        11'd1559: data_font_rom = 8'b01111100; // 7  *****
        11'd1560: data_font_rom = 8'b11001100; // 8 **  **
        11'd1561: data_font_rom = 8'b11001100; // 9 **  **
        11'd1562: data_font_rom = 8'b11001100; // a **  **
        11'd1563: data_font_rom = 8'b01110110; // b  *** **
        11'd1564: data_font_rom = 8'b00000000; // c
        11'd1565: data_font_rom = 8'b00000000; // d
        11'd1566: data_font_rom = 8'b00000000; // e
        11'd1567: data_font_rom = 8'b00000000; // f
        // code x62
        11'd1568: data_font_rom = 8'b00000000; // 0
        11'd1569: data_font_rom = 8'b00000000; // 1
        11'd1570: data_font_rom = 8'b11100000; // 2  ***
        11'd1571: data_font_rom = 8'b01100000; // 3   **
        11'd1572: data_font_rom = 8'b01100000; // 4   **
        11'd1573: data_font_rom = 8'b01111000; // 5   ****
        11'd1574: data_font_rom = 8'b01101100; // 6   ** **
        11'd1575: data_font_rom = 8'b01100110; // 7   **  **
        11'd1576: data_font_rom = 8'b01100110; // 8   **  **
        11'd1577: data_font_rom = 8'b01100110; // 9   **  **
        11'd1578: data_font_rom = 8'b01100110; // a   **  **
        11'd1579: data_font_rom = 8'b01111100; // b   *****
        11'd1580: data_font_rom = 8'b00000000; // c
        11'd1581: data_font_rom = 8'b00000000; // d
        11'd1582: data_font_rom = 8'b00000000; // e
        11'd1583: data_font_rom = 8'b00000000; // f
        // code x63
        11'd1584: data_font_rom = 8'b00000000; // 0
        11'd1585: data_font_rom = 8'b00000000; // 1
        11'd1586: data_font_rom = 8'b00000000; // 2
        11'd1587: data_font_rom = 8'b00000000; // 3
        11'd1588: data_font_rom = 8'b00000000; // 4
        11'd1589: data_font_rom = 8'b01111100; // 5  *****
        11'd1590: data_font_rom = 8'b11000110; // 6 **   **
        11'd1591: data_font_rom = 8'b11000000; // 7 **
        11'd1592: data_font_rom = 8'b11000000; // 8 **
        11'd1593: data_font_rom = 8'b11000000; // 9 **
        11'd1594: data_font_rom = 8'b11000110; // a **   **
        11'd1595: data_font_rom = 8'b01111100; // b  *****
        11'd1596: data_font_rom = 8'b00000000; // c
        11'd1597: data_font_rom = 8'b00000000; // d
        11'd1598: data_font_rom = 8'b00000000; // e
        11'd1599: data_font_rom = 8'b00000000; // f
        // code x64
        11'd1600: data_font_rom = 8'b00000000; // 0
        11'd1601: data_font_rom = 8'b00000000; // 1
        11'd1602: data_font_rom = 8'b00011100; // 2    ***
        11'd1603: data_font_rom = 8'b00001100; // 3     **
        11'd1604: data_font_rom = 8'b00001100; // 4     **
        11'd1605: data_font_rom = 8'b00111100; // 5   ****
        11'd1606: data_font_rom = 8'b01101100; // 6  ** **
        11'd1607: data_font_rom = 8'b11001100; // 7 **  **
        11'd1608: data_font_rom = 8'b11001100; // 8 **  **
        11'd1609: data_font_rom = 8'b11001100; // 9 **  **
        11'd1610: data_font_rom = 8'b11001100; // a **  **
        11'd1611: data_font_rom = 8'b01110110; // b  *** **
        11'd1612: data_font_rom = 8'b00000000; // c
        11'd1613: data_font_rom = 8'b00000000; // d
        11'd1614: data_font_rom = 8'b00000000; // e
        11'd1615: data_font_rom = 8'b00000000; // f
        // code x65
        11'd1616: data_font_rom = 8'b00000000; // 0
        11'd1617: data_font_rom = 8'b00000000; // 1
        11'd1618: data_font_rom = 8'b00000000; // 2
        11'd1619: data_font_rom = 8'b00000000; // 3
        11'd1620: data_font_rom = 8'b00000000; // 4
        11'd1621: data_font_rom = 8'b01111100; // 5  *****
        11'd1622: data_font_rom = 8'b11000110; // 6 **   **
        11'd1623: data_font_rom = 8'b11111110; // 7 *******
        11'd1624: data_font_rom = 8'b11000000; // 8 **
        11'd1625: data_font_rom = 8'b11000000; // 9 **
        11'd1626: data_font_rom = 8'b11000110; // a **   **
        11'd1627: data_font_rom = 8'b01111100; // b  *****
        11'd1628: data_font_rom = 8'b00000000; // c
        11'd1629: data_font_rom = 8'b00000000; // d
        11'd1630: data_font_rom = 8'b00000000; // e
        11'd1631: data_font_rom = 8'b00000000; // f
        // code x66
        11'd1632: data_font_rom = 8'b00000000; // 0
        11'd1633: data_font_rom = 8'b00000000; // 1
        11'd1634: data_font_rom = 8'b00111000; // 2   ***
        11'd1635: data_font_rom = 8'b01101100; // 3  ** **
        11'd1636: data_font_rom = 8'b01100100; // 4  **  *
        11'd1637: data_font_rom = 8'b01100000; // 5  **
        11'd1638: data_font_rom = 8'b11110000; // 6 ****
        11'd1639: data_font_rom = 8'b01100000; // 7  **
        11'd1640: data_font_rom = 8'b01100000; // 8  **
        11'd1641: data_font_rom = 8'b01100000; // 9  **
        11'd1642: data_font_rom = 8'b01100000; // a  **
        11'd1643: data_font_rom = 8'b11110000; // b ****
        11'd1644: data_font_rom = 8'b00000000; // c
        11'd1645: data_font_rom = 8'b00000000; // d
        11'd1646: data_font_rom = 8'b00000000; // e
        11'd1647: data_font_rom = 8'b00000000; // f
        // code x67
        11'd1648: data_font_rom = 8'b00000000; // 0
        11'd1649: data_font_rom = 8'b00000000; // 1
        11'd1650: data_font_rom = 8'b00000000; // 2
        11'd1651: data_font_rom = 8'b00000000; // 3
        11'd1652: data_font_rom = 8'b00000000; // 4
        11'd1653: data_font_rom = 8'b01110110; // 5  *** **
        11'd1654: data_font_rom = 8'b11001100; // 6 **  **
        11'd1655: data_font_rom = 8'b11001100; // 7 **  **
        11'd1656: data_font_rom = 8'b11001100; // 8 **  **
        11'd1657: data_font_rom = 8'b11001100; // 9 **  **
        11'd1658: data_font_rom = 8'b11001100; // a **  **
        11'd1659: data_font_rom = 8'b01111100; // b  *****
        11'd1660: data_font_rom = 8'b00001100; // c     **
        11'd1661: data_font_rom = 8'b11001100; // d **  **
        11'd1662: data_font_rom = 8'b01111000; // e  ****
        11'd1663: data_font_rom = 8'b00000000; // f
        // code x68
        11'd1664: data_font_rom = 8'b00000000; // 0
        11'd1665: data_font_rom = 8'b00000000; // 1
        11'd1666: data_font_rom = 8'b11100000; // 2 ***
        11'd1667: data_font_rom = 8'b01100000; // 3  **
        11'd1668: data_font_rom = 8'b01100000; // 4  **
        11'd1669: data_font_rom = 8'b01101100; // 5  ** **
        11'd1670: data_font_rom = 8'b01110110; // 6  *** **
        11'd1671: data_font_rom = 8'b01100110; // 7  **  **
        11'd1672: data_font_rom = 8'b01100110; // 8  **  **
        11'd1673: data_font_rom = 8'b01100110; // 9  **  **
        11'd1674: data_font_rom = 8'b01100110; // a  **  **
        11'd1675: data_font_rom = 8'b11100110; // b ***  **
        11'd1676: data_font_rom = 8'b00000000; // c
        11'd1677: data_font_rom = 8'b00000000; // d
        11'd1678: data_font_rom = 8'b00000000; // e
        11'd1679: data_font_rom = 8'b00000000; // f
        // code x69
        11'd1680: data_font_rom = 8'b00000000; // 0
        11'd1681: data_font_rom = 8'b00000000; // 1
        11'd1682: data_font_rom = 8'b00011000; // 2    **
        11'd1683: data_font_rom = 8'b00011000; // 3    **
        11'd1684: data_font_rom = 8'b00000000; // 4
        11'd1685: data_font_rom = 8'b00111000; // 5   ***
        11'd1686: data_font_rom = 8'b00011000; // 6    **
        11'd1687: data_font_rom = 8'b00011000; // 7    **
        11'd1688: data_font_rom = 8'b00011000; // 8    **
        11'd1689: data_font_rom = 8'b00011000; // 9    **
        11'd1690: data_font_rom = 8'b00011000; // a    **
        11'd1691: data_font_rom = 8'b00111100; // b   ****
        11'd1692: data_font_rom = 8'b00000000; // c
        11'd1693: data_font_rom = 8'b00000000; // d
        11'd1694: data_font_rom = 8'b00000000; // e
        11'd1695: data_font_rom = 8'b00000000; // f
        // code x6a
        11'd1696: data_font_rom = 8'b00000000; // 0
        11'd1697: data_font_rom = 8'b00000000; // 1
        11'd1698: data_font_rom = 8'b00000110; // 2      **
        11'd1699: data_font_rom = 8'b00000110; // 3      **
        11'd1700: data_font_rom = 8'b00000000; // 4
        11'd1701: data_font_rom = 8'b00001110; // 5     ***
        11'd1702: data_font_rom = 8'b00000110; // 6      **
        11'd1703: data_font_rom = 8'b00000110; // 7      **
        11'd1704: data_font_rom = 8'b00000110; // 8      **
        11'd1705: data_font_rom = 8'b00000110; // 9      **
        11'd1706: data_font_rom = 8'b00000110; // a      **
        11'd1707: data_font_rom = 8'b00000110; // b      **
        11'd1708: data_font_rom = 8'b01100110; // c  **  **
        11'd1709: data_font_rom = 8'b01100110; // d  **  **
        11'd1710: data_font_rom = 8'b00111100; // e   ****
        11'd1711: data_font_rom = 8'b00000000; // f
        // code x6b
        11'd1712: data_font_rom = 8'b00000000; // 0
        11'd1713: data_font_rom = 8'b00000000; // 1
        11'd1714: data_font_rom = 8'b11100000; // 2 ***
        11'd1715: data_font_rom = 8'b01100000; // 3  **
        11'd1716: data_font_rom = 8'b01100000; // 4  **
        11'd1717: data_font_rom = 8'b01100110; // 5  **  **
        11'd1718: data_font_rom = 8'b01101100; // 6  ** **
        11'd1719: data_font_rom = 8'b01111000; // 7  ****
        11'd1720: data_font_rom = 8'b01111000; // 8  ****
        11'd1721: data_font_rom = 8'b01101100; // 9  ** **
        11'd1722: data_font_rom = 8'b01100110; // a  **  **
        11'd1723: data_font_rom = 8'b11100110; // b ***  **
        11'd1724: data_font_rom = 8'b00000000; // c
        11'd1725: data_font_rom = 8'b00000000; // d
        11'd1726: data_font_rom = 8'b00000000; // e
        11'd1727: data_font_rom = 8'b00000000; // f
        // code x6c
        11'd1728: data_font_rom = 8'b00000000; // 0
        11'd1729: data_font_rom = 8'b00000000; // 1
        11'd1730: data_font_rom = 8'b00111000; // 2   ***
        11'd1731: data_font_rom = 8'b00011000; // 3    **
        11'd1732: data_font_rom = 8'b00011000; // 4    **
        11'd1733: data_font_rom = 8'b00011000; // 5    **
        11'd1734: data_font_rom = 8'b00011000; // 6    **
        11'd1735: data_font_rom = 8'b00011000; // 7    **
        11'd1736: data_font_rom = 8'b00011000; // 8    **
        11'd1737: data_font_rom = 8'b00011000; // 9    **
        11'd1738: data_font_rom = 8'b00011000; // a    **
        11'd1739: data_font_rom = 8'b00111100; // b   ****
        11'd1740: data_font_rom = 8'b00000000; // c
        11'd1741: data_font_rom = 8'b00000000; // d
        11'd1742: data_font_rom = 8'b00000000; // e
        11'd1743: data_font_rom = 8'b00000000; // f
        // code x6d
        11'd1744: data_font_rom = 8'b00000000; // 0
        11'd1745: data_font_rom = 8'b00000000; // 1
        11'd1746: data_font_rom = 8'b00000000; // 2
        11'd1747: data_font_rom = 8'b00000000; // 3
        11'd1748: data_font_rom = 8'b00000000; // 4
        11'd1749: data_font_rom = 8'b11100110; // 5 ***  **
        11'd1750: data_font_rom = 8'b11111111; // 6 ********
        11'd1751: data_font_rom = 8'b11011011; // 7 ** ** **
        11'd1752: data_font_rom = 8'b11011011; // 8 ** ** **
        11'd1753: data_font_rom = 8'b11011011; // 9 ** ** **
        11'd1754: data_font_rom = 8'b11011011; // a ** ** **
        11'd1755: data_font_rom = 8'b11011011; // b ** ** **
        11'd1756: data_font_rom = 8'b00000000; // c
        11'd1757: data_font_rom = 8'b00000000; // d
        11'd1758: data_font_rom = 8'b00000000; // e
        11'd1759: data_font_rom = 8'b00000000; // f
        // code x6e
        11'd1760: data_font_rom = 8'b00000000; // 0
        11'd1761: data_font_rom = 8'b00000000; // 1
        11'd1762: data_font_rom = 8'b00000000; // 2
        11'd1763: data_font_rom = 8'b00000000; // 3
        11'd1764: data_font_rom = 8'b00000000; // 4
        11'd1765: data_font_rom = 8'b11011100; // 5 ** ***
        11'd1766: data_font_rom = 8'b01100110; // 6  **  **
        11'd1767: data_font_rom = 8'b01100110; // 7  **  **
        11'd1768: data_font_rom = 8'b01100110; // 8  **  **
        11'd1769: data_font_rom = 8'b01100110; // 9  **  **
        11'd1770: data_font_rom = 8'b01100110; // a  **  **
        11'd1771: data_font_rom = 8'b01100110; // b  **  **
        11'd1772: data_font_rom = 8'b00000000; // c
        11'd1773: data_font_rom = 8'b00000000; // d
        11'd1774: data_font_rom = 8'b00000000; // e
        11'd1775: data_font_rom = 8'b00000000; // f
        // code x6f
        11'd1776: data_font_rom = 8'b00000000; // 0
        11'd1777: data_font_rom = 8'b00000000; // 1
        11'd1778: data_font_rom = 8'b00000000; // 2
        11'd1779: data_font_rom = 8'b00000000; // 3
        11'd1780: data_font_rom = 8'b00000000; // 4
        11'd1781: data_font_rom = 8'b01111100; // 5  *****
        11'd1782: data_font_rom = 8'b11000110; // 6 **   **
        11'd1783: data_font_rom = 8'b11000110; // 7 **   **
        11'd1784: data_font_rom = 8'b11000110; // 8 **   **
        11'd1785: data_font_rom = 8'b11000110; // 9 **   **
        11'd1786: data_font_rom = 8'b11000110; // a **   **
        11'd1787: data_font_rom = 8'b01111100; // b  *****
        11'd1788: data_font_rom = 8'b00000000; // c
        11'd1789: data_font_rom = 8'b00000000; // d
        11'd1790: data_font_rom = 8'b00000000; // e
        11'd1791: data_font_rom = 8'b00000000; // f
        // code x70
        11'd1792: data_font_rom = 8'b00000000; // 0
        11'd1793: data_font_rom = 8'b00000000; // 1
        11'd1794: data_font_rom = 8'b00000000; // 2
        11'd1795: data_font_rom = 8'b00000000; // 3
        11'd1796: data_font_rom = 8'b00000000; // 4
        11'd1797: data_font_rom = 8'b11011100; // 5 ** ***
        11'd1798: data_font_rom = 8'b01100110; // 6  **  **
        11'd1799: data_font_rom = 8'b01100110; // 7  **  **
        11'd1800: data_font_rom = 8'b01100110; // 8  **  **
        11'd1801: data_font_rom = 8'b01100110; // 9  **  **
        11'd1802: data_font_rom = 8'b01100110; // a  **  **
        11'd1803: data_font_rom = 8'b01111100; // b  *****
        11'd1804: data_font_rom = 8'b01100000; // c  **
        11'd1805: data_font_rom = 8'b01100000; // d  **
        11'd1806: data_font_rom = 8'b11110000; // e ****
        11'd1807: data_font_rom = 8'b00000000; // f
        // code x71
        11'd1808: data_font_rom = 8'b00000000; // 0
        11'd1809: data_font_rom = 8'b00000000; // 1
        11'd1810: data_font_rom = 8'b00000000; // 2
        11'd1811: data_font_rom = 8'b00000000; // 3
        11'd1812: data_font_rom = 8'b00000000; // 4
        11'd1813: data_font_rom = 8'b01110110; // 5  *** **
        11'd1814: data_font_rom = 8'b11001100; // 6 **  **
        11'd1815: data_font_rom = 8'b11001100; // 7 **  **
        11'd1816: data_font_rom = 8'b11001100; // 8 **  **
        11'd1817: data_font_rom = 8'b11001100; // 9 **  **
        11'd1818: data_font_rom = 8'b11001100; // a **  **
        11'd1819: data_font_rom = 8'b01111100; // b  *****
        11'd1820: data_font_rom = 8'b00001100; // c     **
        11'd1821: data_font_rom = 8'b00001100; // d     **
        11'd1822: data_font_rom = 8'b00011110; // e    ****
        11'd1823: data_font_rom = 8'b00000000; // f
        // code x72
        11'd1824: data_font_rom = 8'b00000000; // 0
        11'd1825: data_font_rom = 8'b00000000; // 1
        11'd1826: data_font_rom = 8'b00000000; // 2
        11'd1827: data_font_rom = 8'b00000000; // 3
        11'd1828: data_font_rom = 8'b00000000; // 4
        11'd1829: data_font_rom = 8'b11011100; // 5 ** ***
        11'd1830: data_font_rom = 8'b01110110; // 6  *** **
        11'd1831: data_font_rom = 8'b01100110; // 7  **  **
        11'd1832: data_font_rom = 8'b01100000; // 8  **
        11'd1833: data_font_rom = 8'b01100000; // 9  **
        11'd1834: data_font_rom = 8'b01100000; // a  **
        11'd1835: data_font_rom = 8'b11110000; // b ****
        11'd1836: data_font_rom = 8'b00000000; // c
        11'd1837: data_font_rom = 8'b00000000; // d
        11'd1838: data_font_rom = 8'b00000000; // e
        11'd1839: data_font_rom = 8'b00000000; // f
        // code x73
        11'd1840: data_font_rom = 8'b00000000; // 0
        11'd1841: data_font_rom = 8'b00000000; // 1
        11'd1842: data_font_rom = 8'b00000000; // 2
        11'd1843: data_font_rom = 8'b00000000; // 3
        11'd1844: data_font_rom = 8'b00000000; // 4
        11'd1845: data_font_rom = 8'b01111100; // 5  *****
        11'd1846: data_font_rom = 8'b11000110; // 6 **   **
        11'd1847: data_font_rom = 8'b01100000; // 7  **
        11'd1848: data_font_rom = 8'b00111000; // 8   ***
        11'd1849: data_font_rom = 8'b00001100; // 9     **
        11'd1850: data_font_rom = 8'b11000110; // a **   **
        11'd1851: data_font_rom = 8'b01111100; // b  *****
        11'd1852: data_font_rom = 8'b00000000; // c
        11'd1853: data_font_rom = 8'b00000000; // d
        11'd1854: data_font_rom = 8'b00000000; // e
        11'd1855: data_font_rom = 8'b00000000; // f
        // code x74
        11'd1856: data_font_rom = 8'b00000000; // 0
        11'd1857: data_font_rom = 8'b00000000; // 1
        11'd1858: data_font_rom = 8'b00010000; // 2    *
        11'd1859: data_font_rom = 8'b00110000; // 3   **
        11'd1860: data_font_rom = 8'b00110000; // 4   **
        11'd1861: data_font_rom = 8'b11111100; // 5 ******
        11'd1862: data_font_rom = 8'b00110000; // 6   **
        11'd1863: data_font_rom = 8'b00110000; // 7   **
        11'd1864: data_font_rom = 8'b00110000; // 8   **
        11'd1865: data_font_rom = 8'b00110000; // 9   **
        11'd1866: data_font_rom = 8'b00110110; // a   ** **
        11'd1867: data_font_rom = 8'b00011100; // b    ***
        11'd1868: data_font_rom = 8'b00000000; // c
        11'd1869: data_font_rom = 8'b00000000; // d
        11'd1870: data_font_rom = 8'b00000000; // e
        11'd1871: data_font_rom = 8'b00000000; // f
        // code x75
        11'd1872: data_font_rom = 8'b00000000; // 0
        11'd1873: data_font_rom = 8'b00000000; // 1
        11'd1874: data_font_rom = 8'b00000000; // 2
        11'd1875: data_font_rom = 8'b00000000; // 3
        11'd1876: data_font_rom = 8'b00000000; // 4
        11'd1877: data_font_rom = 8'b11001100; // 5 **  **
        11'd1878: data_font_rom = 8'b11001100; // 6 **  **
        11'd1879: data_font_rom = 8'b11001100; // 7 **  **
        11'd1880: data_font_rom = 8'b11001100; // 8 **  **
        11'd1881: data_font_rom = 8'b11001100; // 9 **  **
        11'd1882: data_font_rom = 8'b11001100; // a **  **
        11'd1883: data_font_rom = 8'b01110110; // b  *** **
        11'd1884: data_font_rom = 8'b00000000; // c
        11'd1885: data_font_rom = 8'b00000000; // d
        11'd1886: data_font_rom = 8'b00000000; // e
        11'd1887: data_font_rom = 8'b00000000; // f
        // code x76
        11'd1888: data_font_rom = 8'b00000000; // 0
        11'd1889: data_font_rom = 8'b00000000; // 1
        11'd1890: data_font_rom = 8'b00000000; // 2
        11'd1891: data_font_rom = 8'b00000000; // 3
        11'd1892: data_font_rom = 8'b00000000; // 4
        11'd1893: data_font_rom = 8'b11000011; // 5 **    **
        11'd1894: data_font_rom = 8'b11000011; // 6 **    **
        11'd1895: data_font_rom = 8'b11000011; // 7 **    **
        11'd1896: data_font_rom = 8'b11000011; // 8 **    **
        11'd1897: data_font_rom = 8'b01100110; // 9  **  **
        11'd1898: data_font_rom = 8'b00111100; // a   ****
        11'd1899: data_font_rom = 8'b00011000; // b    **
        11'd1900: data_font_rom = 8'b00000000; // c
        11'd1901: data_font_rom = 8'b00000000; // d
        11'd1902: data_font_rom = 8'b00000000; // e
        11'd1903: data_font_rom = 8'b00000000; // f
        // code x77
        11'd1904: data_font_rom = 8'b00000000; // 0
        11'd1905: data_font_rom = 8'b00000000; // 1
        11'd1906: data_font_rom = 8'b00000000; // 2
        11'd1907: data_font_rom = 8'b00000000; // 3
        11'd1908: data_font_rom = 8'b00000000; // 4
        11'd1909: data_font_rom = 8'b11000011; // 5 **    **
        11'd1910: data_font_rom = 8'b11000011; // 6 **    **
        11'd1911: data_font_rom = 8'b11000011; // 7 **    **
        11'd1912: data_font_rom = 8'b11011011; // 8 ** ** **
        11'd1913: data_font_rom = 8'b11011011; // 9 ** ** **
        11'd1914: data_font_rom = 8'b11111111; // a ********
        11'd1915: data_font_rom = 8'b01100110; // b  **  **
        11'd1916: data_font_rom = 8'b00000000; // c
        11'd1917: data_font_rom = 8'b00000000; // d
        11'd1918: data_font_rom = 8'b00000000; // e
        11'd1919: data_font_rom = 8'b00000000; // f
        // code x78
        11'd1920: data_font_rom = 8'b00000000; // 0
        11'd1921: data_font_rom = 8'b00000000; // 1
        11'd1922: data_font_rom = 8'b00000000; // 2
        11'd1923: data_font_rom = 8'b00000000; // 3
        11'd1924: data_font_rom = 8'b00000000; // 4
        11'd1925: data_font_rom = 8'b11000011; // 5 **    **
        11'd1926: data_font_rom = 8'b01100110; // 6  **  **
        11'd1927: data_font_rom = 8'b00111100; // 7   ****
        11'd1928: data_font_rom = 8'b00011000; // 8    **
        11'd1929: data_font_rom = 8'b00111100; // 9   ****
        11'd1930: data_font_rom = 8'b01100110; // a  **  **
        11'd1931: data_font_rom = 8'b11000011; // b **    **
        11'd1932: data_font_rom = 8'b00000000; // c
        11'd1933: data_font_rom = 8'b00000000; // d
        11'd1934: data_font_rom = 8'b00000000; // e
        11'd1935: data_font_rom = 8'b00000000; // f
        // code x79
        11'd1936: data_font_rom = 8'b00000000; // 0
        11'd1937: data_font_rom = 8'b00000000; // 1
        11'd1938: data_font_rom = 8'b00000000; // 2
        11'd1939: data_font_rom = 8'b00000000; // 3
        11'd1940: data_font_rom = 8'b00000000; // 4
        11'd1941: data_font_rom = 8'b11000110; // 5 **   **
        11'd1942: data_font_rom = 8'b11000110; // 6 **   **
        11'd1943: data_font_rom = 8'b11000110; // 7 **   **
        11'd1944: data_font_rom = 8'b11000110; // 8 **   **
        11'd1945: data_font_rom = 8'b11000110; // 9 **   **
        11'd1946: data_font_rom = 8'b11000110; // a **   **
        11'd1947: data_font_rom = 8'b01111110; // b  ******
        11'd1948: data_font_rom = 8'b00000110; // c      **
        11'd1949: data_font_rom = 8'b00001100; // d     **
        11'd1950: data_font_rom = 8'b11111000; // e *****
        11'd1951: data_font_rom = 8'b00000000; // f
        // code x7a
        11'd1952: data_font_rom = 8'b00000000; // 0
        11'd1953: data_font_rom = 8'b00000000; // 1
        11'd1954: data_font_rom = 8'b00000000; // 2
        11'd1955: data_font_rom = 8'b00000000; // 3
        11'd1956: data_font_rom = 8'b00000000; // 4
        11'd1957: data_font_rom = 8'b11111110; // 5 *******
        11'd1958: data_font_rom = 8'b11001100; // 6 **  **
        11'd1959: data_font_rom = 8'b00011000; // 7    **
        11'd1960: data_font_rom = 8'b00110000; // 8   **
        11'd1961: data_font_rom = 8'b01100000; // 9  **
        11'd1962: data_font_rom = 8'b11000110; // a **   **
        11'd1963: data_font_rom = 8'b11111110; // b *******
        11'd1964: data_font_rom = 8'b00000000; // c
        11'd1965: data_font_rom = 8'b00000000; // d
        11'd1966: data_font_rom = 8'b00000000; // e
        11'd1967: data_font_rom = 8'b00000000; // f
        // code x7b
        11'd1968: data_font_rom = 8'b00000000; // 0
        11'd1969: data_font_rom = 8'b00000000; // 1
        11'd1970: data_font_rom = 8'b00001110; // 2     ***
        11'd1971: data_font_rom = 8'b00011000; // 3    **
        11'd1972: data_font_rom = 8'b00011000; // 4    **
        11'd1973: data_font_rom = 8'b00011000; // 5    **
        11'd1974: data_font_rom = 8'b01110000; // 6  ***
        11'd1975: data_font_rom = 8'b00011000; // 7    **
        11'd1976: data_font_rom = 8'b00011000; // 8    **
        11'd1977: data_font_rom = 8'b00011000; // 9    **
        11'd1978: data_font_rom = 8'b00011000; // a    **
        11'd1979: data_font_rom = 8'b00001110; // b     ***
        11'd1980: data_font_rom = 8'b00000000; // c
        11'd1981: data_font_rom = 8'b00000000; // d
        11'd1982: data_font_rom = 8'b00000000; // e
        11'd1983: data_font_rom = 8'b00000000; // f
        // code x7c
        11'd1984: data_font_rom = 8'b00000000; // 0
        11'd1985: data_font_rom = 8'b00000000; // 1
        11'd1986: data_font_rom = 8'b00011000; // 2    **
        11'd1987: data_font_rom = 8'b00011000; // 3    **
        11'd1988: data_font_rom = 8'b00011000; // 4    **
        11'd1989: data_font_rom = 8'b00011000; // 5    **
        11'd1990: data_font_rom = 8'b00000000; // 6
        11'd1991: data_font_rom = 8'b00011000; // 7    **
        11'd1992: data_font_rom = 8'b00011000; // 8    **
        11'd1993: data_font_rom = 8'b00011000; // 9    **
        11'd1994: data_font_rom = 8'b00011000; // a    **
        11'd1995: data_font_rom = 8'b00011000; // b    **
        11'd1996: data_font_rom = 8'b00000000; // c
        11'd1997: data_font_rom = 8'b00000000; // d
        11'd1998: data_font_rom = 8'b00000000; // e
        11'd1999: data_font_rom = 8'b00000000; // f
        // code x7d
        11'd2000: data_font_rom = 8'b00000000; // 0
        11'd2001: data_font_rom = 8'b00000000; // 1
        11'd2002: data_font_rom = 8'b01110000; // 2  ***
        11'd2003: data_font_rom = 8'b00011000; // 3    **
        11'd2004: data_font_rom = 8'b00011000; // 4    **
        11'd2005: data_font_rom = 8'b00011000; // 5    **
        11'd2006: data_font_rom = 8'b00001110; // 6     ***
        11'd2007: data_font_rom = 8'b00011000; // 7    **
        11'd2008: data_font_rom = 8'b00011000; // 8    **
        11'd2009: data_font_rom = 8'b00011000; // 9    **
        11'd2010: data_font_rom = 8'b00011000; // a    **
        11'd2011: data_font_rom = 8'b01110000; // b  ***
        11'd2012: data_font_rom = 8'b00000000; // c
        11'd2013: data_font_rom = 8'b00000000; // d
        11'd2014: data_font_rom = 8'b00000000; // e
        11'd2015: data_font_rom = 8'b00000000; // f
        // code x7e
        11'd2016: data_font_rom = 8'b00000000; // 0
        11'd2017: data_font_rom = 8'b00000000; // 1
        11'd2018: data_font_rom = 8'b01110110; // 2  *** **
        11'd2019: data_font_rom = 8'b11011100; // 3 ** ***
        11'd2020: data_font_rom = 8'b00000000; // 4
        11'd2021: data_font_rom = 8'b00000000; // 5
        11'd2022: data_font_rom = 8'b00000000; // 6
        11'd2023: data_font_rom = 8'b00000000; // 7
        11'd2024: data_font_rom = 8'b00000000; // 8
        11'd2025: data_font_rom = 8'b00000000; // 9
        11'd2026: data_font_rom = 8'b00000000; // a
        11'd2027: data_font_rom = 8'b00000000; // b
        11'd2028: data_font_rom = 8'b00000000; // c
        11'd2029: data_font_rom = 8'b00000000; // d
        11'd2030: data_font_rom = 8'b00000000; // e
        11'd2031: data_font_rom = 8'b00000000; // f
        // code x7f
        11'd2032: data_font_rom = 8'b00000000; // 0
        11'd2033: data_font_rom = 8'b00000000; // 1
        11'd2034: data_font_rom = 8'b00000000; // 2
        11'd2035: data_font_rom = 8'b00000000; // 3
        11'd2036: data_font_rom = 8'b00010000; // 4    *
        11'd2037: data_font_rom = 8'b00111000; // 5   ***
        11'd2038: data_font_rom = 8'b01101100; // 6  ** **
        11'd2039: data_font_rom = 8'b11000110; // 7 **   **
        11'd2040: data_font_rom = 8'b11000110; // 8 **   **
        11'd2041: data_font_rom = 8'b11000110; // 9 **   **
        11'd2042: data_font_rom = 8'b11111110; // a *******
        11'd2043: data_font_rom = 8'b00000000; // b
        11'd2044: data_font_rom = 8'b00000000; // c
        11'd2045: data_font_rom = 8'b00000000; // d
        11'd2046: data_font_rom = 8'b00000000; // e
        11'd2047: data_font_rom = 8'b00000000;  // f
    endcase

endmodule
